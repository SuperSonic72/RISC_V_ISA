----------------------------------------------------------------------------------
-- Company: Covnetics Limited (at the time of development)
-- Engineer: ED72
-- 
-- Create Date:    09:33:24 18/10/2022 
-- Design Name: 
-- Module Name:    RISC_V_Core - Behavioral 
-- Project Name:   RISC_V
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--
--
entity RISC_V_Core is
    Port ( RST           : in  std_logic;                       -- Reset signal
           CLK           : in  std_logic;                       -- Clock signal
           CONTR_OUT     : out std_logic_vector(31 downto 0);   -- Control Output - used in validation
           PORT_A        : out std_logic_vector(31 downto 0)    -- Processor general purpose port - Memory mapped at 0x0000
     );
end RISC_V_Core;
--
--
architecture Behavioral of RISC_V_Core is
--
	  -- Enumerated operation
	  type RISC_V_OPERATION is 
	  (o_SUM, o_SUB, o_SHIFT_LEFT, o_SHIFT_RIGHT, o_SRA, o_AND, o_OR, o_XOR, o_SLT, o_SLTU, o_LOAD, o_SAVE);
	  type DATA_F is 
	  (l_32, l_16, l_8, l_16_U, l_8_U);
--
	  type X_REG is array (0 to 31) of signed(31 downto 0);
	  type RAM_MEM_1 is array (0 to 2047) of std_logic_vector(31 downto 0);
	  type RAM_MEM_2 is array (0 to 1023) of std_logic_vector(31 downto 0);
--
	  signal   OPERATION             : RISC_V_OPERATION;
      signal   PROG_MEM              : RAM_MEM_1 := 
(X"740A4661",X"6D696C79",X"3A205472",X"696F6E0A",X"44657669",X"63653A20",X"54384638",X"310A5769",X"6474683A",X"20310A50",X"41444445",
X"445F4249",X"54533A20",X"300A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",
X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",
X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"168A2236",X"FFFE0740",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00010000",X"00000001",
X"00000000",X"00000000",X"00358341",X"50100060",X"00152200",X"002AC855",X"90AB2156",X"42AC8559",X"08311564",X"2AC85590",X"AB215642",
X"AC85590A",X"B2106220",X"4C559083",X"1106220C",X"44188831",X"10622AC8",X"5590AB21",X"5642AC85",X"590AB215",X"642AC851",X"90813146",
X"429CB002",X"60E4F041",X"88A32156",X"420C4559",X"0AB21564",X"2AC85590",X"AB215642",X"AC84098A",X"B2156420",X"A0559082",X"81026206",
X"C40D8AB2",X"00000000",X"00000000",X"00000000",X"90088082",X"40A09048",X"04122800",X"82410090",X"48241201",X"048A4120",X"00090480",
X"41209049",X"64120904",X"82492090",X"48241209",X"04824122",X"00090482",X"41209020",X"24060904",X"82410090",X"08240605",X"01920922",
X"90090482",X"41021248",X"240A7114",X"88406290",X"48A41229",X"04924122",X"9009048A",X"41239049",X"14500824",X"96412080",X"48241209",
X"04020120",X"00090480",X"41229048",X"24120904",X"82412090",X"48044209",X"148A4B20",X"00090482",X"41209148",X"0C920904",X"82412090",
X"48240221",X"04824520",X"90090482",X"41209048",X"20120134",X"82112590",X"48041209",X"00824100",X"00000000",X"00000000",X"00000000",
X"00001000",X"00000000",X"10000102",X"00081000",X"00000002",X"00140000",X"00000000",X"80000000",X"80000000",X"00040000",X"00000000",
X"00000001",X"00000000",X"00000004",X"00000000",X"00002000",X"10000000",X"00081401",X"00000000",X"08140100",X"00006220",X"10000700",
X"00000050",X"001C0001",X"00000004",X"00070000",X"80820110",X"080A0008",X"00000000",X"00801005",X"00000010",X"80040000",X"00000000",
X"00000000",X"00088800",X"00100400",X"00000000",X"00000000",X"00400000",X"00000000",X"00000440",X"00000000",X"00000000",X"00000000",
X"04000210",X"00000000",X"00200000",X"01000010",X"00000000",X"00000000",X"00000000",X"90093490",X"49248209",X"24B2092C",X"92492592",
X"C9E41209",X"14824121",X"00092482",X"49259048",X"24120904",X"80412090",X"48241209",X"04824125",X"00090482",X"41209049",X"C4B23824",
X"12412190",X"49224249",X"34820B20",X"90090496",X"41020148",X"0C824824",X"82052612",X"48248229",X"00024124",X"90082482",X"49209018",
X"1450432C",X"15052092",X"C8241079",X"048A4F20",X"00432482",X"45109048",X"04520904",X"924AA290",X"48241209",X"00924120",X"0009044A",
X"41209028",X"A492092A",X"82412090",X"49441271",X"241E4920",X"90090482",X"41209248",X"2490A82C",X"824B0090",X"C8245209",X"041A4B26",
X"00000000",X"00000000",X"00000000",X"0000100A",X"04020540",X"80002000",X"08000001",X"00800000",X"00000002",X"00000000",X"04020000",
X"00000000",X"02000000",X"00000000",X"00000002",X"00000000",X"00000000",X"00402110",X"48000200",X"00000420",X"00004000",X"00000000",
X"00042000",X"00402110",X"00000281",X"00000000",X"04200002",X"00005000",X"04040000",X"00022000",X"08400000",X"00000220",X"00000000",
X"00501000",X"00000000",X"10000000",X"00000000",X"00000000",X"00080000",X"00000000",X"00000200",X"00400010",X"00000000",X"00A00022",
X"10480000",X"00000000",X"00000000",X"00400100",X"00002001",X"00000020",X"00080002",X"00000000",X"00000000",X"00000000",X"00008000",
X"00000000",X"00000008",X"00000100",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000100",X"08402000",X"00000200",X"00800000",X"10000000",X"00000004",X"000A0101",X"00040000",X"000C0000",X"00000400",
X"00020000",X"00000000",X"01090000",X"00804008",X"08000000",X"80000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000400",
X"00004040",X"01000400",X"00000000",X"00020100",X"00400010",X"08000000",X"00000020",X"40000000",X"00000000",X"00000000",X"00200000",
X"00000000",X"00000000",X"00000C00",X"00000000",X"00000000",X"00000000",X"00000000",X"00000100",X"00000000",X"00000000",X"00800000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00050200",X"00204000",X"14000400",
X"010000D0",X"48000000",X"00000000",X"000C0580",X"00800000",X"000C0200",X"00000000",X"20080000",X"00001000",X"00080200",X"00002000",
X"100C0000",X"0000A000",X"20000000",X"00000000",X"00000200",X"01000000",X"00000000",X"02012000",X"00080800",X"00000000",X"000D0480",
X"00A00028",X"34000000",X"00018050",X"40000000",X"00000000",X"00040200",X"00800000",X"10000000",X"00000000",X"00080200",X"00000000",
X"00000000",X"00000000",X"048CC86C",X"92190C92",X"41209068",X"64120D04",X"A2412094",X"48241209",X"00004824",X"32090482",X"41209048",
X"24120904",X"82412090",X"48241209",X"00004824",X"120944A3",X"41A890C8",X"64138904",X"A2512194",X"68643A09",X"04804834",X"12A95F83",
X"493594CD",X"25769924",X"82413090",X"48741219",X"0480C824",X"32090482",X"6B21906A",X"A59A0906",X"82412890",X"4E271A0D",X"00024825",
X"12890482",X"59209048",X"241A0904",X"90188090",X"4A251209",X"00004A24",X"12400242",X"43209049",X"24120904",X"80012800",X"5A241209",
X"04804824",X"12090482",X"432890C8",X"241A0904",X"82512090",X"4AE41389",X"00000000",X"00000000",X"00000000",X"0008C080",X"6022000C",
X"08C00200",X"88004000",X"00000008",X"10000000",X"00000000",X"40000000",X"00000000",X"00600000",X"00000000",X"00000000",X"00000000",
X"00000050",X"00902000",X"00000000",X"4000020A",X"60888000",X"00000100",X"00003610",X"06122814",X"02042018",X"00001000",X"00100020",
X"00000000",X"0008000C",X"24450380",X"00080020",X"00000000",X"0000804C",X"00018002",X"04000000",X"00000000",X"00803000",X"0269A460",
X"00C00000",X"00000000",X"000926C0",X"04000000",X"00000000",X"024010B1",X"90000000",X"00000000",X"00000000",X"02000230",X"00804000",
X"00200000",X"04088030",X"00000000",X"00000000",X"00000000",X"9001201C",X"0F209148",X"0172082C",X"00C40700",X"49845214",X"11814122",
X"0000008A",X"45008110",X"20625824",X"88C10820",X"48A41229",X"00164100",X"0004820A",X"41208500",X"89457100",X"8E042284",X"42240604",
X"081CC412",X"90091002",X"01029049",X"A4404912",X"080F2031",X"4880E401",X"10021122",X"9008101E",X"44229140",X"C048203A",X"000A2591",
X"4420A089",X"04000520",X"0002041E",X"01229008",X"94522911",X"94490290",X"49241200",X"04800F02",X"00025080",X"C4229110",X"01122404",
X"16212080",X"20219279",X"18084060",X"90090482",X"41208848",X"84420904",X"80152090",X"01404600",X"00281000",X"00000000",X"00000000",
X"00000000",X"00083850",X"4A000080",X"08C00100",X"40022000",X"00888021",X"00000004",X"00032C10",X"00100A88",X"01642010",X"040A0008",
X"00000050",X"00980010",X"00000040",X"00000242",X"40A04221",X"0C280001",X"00000000",X"90000084",X"00002180",X"4A110000",X"C0055020",
X"50480000",X"80D08252",X"09880004",X"0000A140",X"0C010209",X"E4E10908",X"20C00402",X"0101B050",X"20421000",X"00002898",X"40040011",
X"00A00028",X"00042400",X"00800003",X"0000AA10",X"00002900",X"08800208",X"00005080",X"20000010",X"01404000",X"31148000",X"00002800",
X"00000000",X"20100000",X"00880000",X"40A40004",X"21008510",X"00000000",X"00000000",X"00000000",X"90089282",X"11209048",X"04320284",
X"84000630",X"28245201",X"01824006",X"00030202",X"41209021",X"88A0050C",X"84004810",X"0964B259",X"04824205",X"00000402",X"41201009",
X"44A65810",X"824A0D02",X"0024A0E8",X"40964100",X"84003014",X"42093042",X"A2080900",X"984A4532",X"08240449",X"08324900",X"90010092",
X"4B250389",X"60D20069",X"4000A041",X"49101203",X"24824085",X"00003438",X"0B208349",X"92120902",X"824C2490",X"08041208",X"04840120",
X"00052C80",X"49161000",X"040A0829",X"82412090",X"0920A051",X"24124884",X"84002482",X"412092A9",X"24C64322",X"92486490",X"41500A41",
X"34148005",X"00000000",X"00000000",X"00000000",X"00002000",X"00000000",X"00400000",X"08210600",X"81000008",X"00080096",X"00000080",
X"00000005",X"84020018",X"08240080",X"10804020",X"00000480",X"00000020",X"00000220",X"904020A0",X"00040030",X"08004860",X"000C0410",
X"0000322A",X"05020000",X"00020004",X"10001001",X"00002080",X"11000C20",X"00040408",X"00001320",X"02C00810",X"0A000012",X"00010000",
X"1000000A",X"00049818",X"04001300",X"80000000",X"08008200",X"40200000",X"80082000",X"00000002",X"04068044",X"10000090",X"00000000",
X"20C09100",X"10840010",X"00088000",X"00000000",X"80402010",X"080C0200",X"00400020",X"188020A0",X"00000000",X"00000000",X"00000000",
X"0001C0E6",X"44201008",X"3F420540",X"8FE5A1DC",X"88C4420D",X"16C84420",X"000DC0C8",X"402110CC",X"261EADC8",X"82F0ABD1",X"88840201",
X"10E845B9",X"00075488",X"40203008",X"37320111",X"E841E3D5",X"FE8403A5",X"CBEC45A0",X"040304E3",X"75B91008",X"045B9106",X"EAE2B810",
X"18173301",X"04804422",X"000DD6A6",X"6038306E",X"A43BBDD4",X"8B71A810",X"08264381",X"008471BA",X"000DC888",X"D0221008",X"37020106",
X"E0402010",X"0804022D",X"C083E020",X"000DC088",X"4020106E",X"84622DC6",X"E3702011",X"6E554A83",X"06EC4538",X"040DC080",X"4020DC08",
X"04022100",X"80422011",X"4C664203",X"18C45031",X"00000000",X"00000000",X"00000000",X"028CC00A",X"0E000000",X"00200000",X"10238200",
X"01008000",X"08440800",X"000C0644",X"080002A7",X"40901CC0",X"02000102",X"81008000",X"30640802",X"0004741C",X"0A050060",X"B3D06020",
X"640B87C1",X"E6400190",X"80540800",X"0000147B",X"33980280",X"0099C014",X"46201500",X"0153E070",X"04000800",X"028C8E3F",X"3C180066",
X"611994CC",X"0F358D00",X"0033D980",X"0000308B",X"0000C014",X"04070000",X"23000006",X"00000000",X"0000006C",X"E8032000",X"00047810",
X"00000027",X"03804446",X"633A0002",X"66915980",X"16740B98",X"00044000",X"0000CC00",X"00004000",X"00000003",X"4480C00C",X"E2623098",
X"00000000",X"00000000",X"00000000",X"0480C06B",X"14000000",X"38000CC0",X"03A062C1",X"1000000C",X"C7400000",X"00020140",X"00000010",
X"2A1C8000",X"02B1D8E0",X"00000000",X"006801B8",X"000F4660",X"00002050",X"031D8001",X"6000CAC8",X"76000584",X"43680190",X"44830663",
X"31502000",X"00058003",X"23A49800",X"10131D00",X"06600000",X"048CC702",X"201A2010",X"00000CC5",X"02F1CA20",X"00221982",X"000331D8",
X"0008C000",X"D0000000",X"3B000006",X"60044000",X"10000004",X"C003B000",X"000CC000",X"80000066",X"334004C1",X"03000000",X"36150882",
X"02600158",X"448CC000",X"00000010",X"00000201",X"00004000",X"0C0C0402",X"02202158",X"00000000",X"00000000",X"00000000",X"000CD6E7",
X"10000000",X"300009A0",X"802998E2",X"000C2000",X"C0540E00",X"000C06C4",X"00241233",X"33102220",X"020910EF",X"00000001",X"08F043BD",
X"000E7518",X"00002035",X"9B803218",X"70408CC0",X"260001E2",X"20D00F74",X"00000578",X"00440209",X"443BD109",X"07201203",X"811FD820",
X"2D184221",X"000DC603",X"30182001",X"09C07CC6",X"63318C20",X"093719A0",X"0093BCCC",X"0002F082",X"AC250000",X"6B800006",X"00002000",
X"00008216",X"F0036C24",X"000C5004",X"06070215",X"BB800667",X"73880010",X"6F111DC1",X"0B780FDE",X"00056800",X"00000010",X"08003200",
X"10020010",X"C038C07F",X"F669BD1A",X"00000000",X"00000000",X"00000000",X"90009036",X"04229000",X"20048904",X"80004010",X"12640561",
X"0C880802",X"0008148A",X"40409288",X"88007200",X"8A4C8D93",X"08840621",X"10284000",X"00005480",X"80228804",X"A0423900",X"200B0C09",
X"2982E070",X"91002825",X"9100148A",X"15220900",X"01042910",X"8940062B",X"10247050",X"502214A0",X"9001149E",X"04220001",X"60C00801",
X"1A401213",X"00A04201",X"11084122",X"00046988",X"45002148",X"91A06900",X"96051090",X"48240508",X"30584024",X"00086488",X"0F240401",
X"41022424",X"81412601",X"081150E5",X"14801A0C",X"91080118",X"11208240",X"04F04114",X"10482620",X"40010049",X"28000427",X"00000000",
X"00000000",X"00000000",X"00082108",X"2A410010",X"04800000",X"001A1482",X"80800024",X"10001424",X"00002810",X"00050141",X"00042101",
X"10040002",X"91100012",X"24020100",X"00020000",X"40450021",X"00806004",X"014E0200",X"81D0C868",X"20010507",X"00006014",X"00048244",
X"20A24001",X"10000E01",X"0000C088",X"0A000005",X"00020008",X"00443048",X"82D20040",X"1C008403",X"03048000",X"08960004",X"00000006",
X"20A24001",X"10000E01",X"0000C088",X"0A000005",X"00020008",X"00443048",X"82D20040",X"1C008403",X"03048000",X"08960004",X"08960004",
X"20A24001",X"10000E01",X"0000C088",X"0A000005",X"00020008",X"00443048",X"82D20040",X"1C008403",X"03048000",X"08960004",X"08960004",
X"00100680",X"00C62001",X"10180000",X"00000001",X"1C0A0102",X"00003814",X"CC022048",X"00844040",X"00000104",X"10008020",X"08960004",X"08960004",
X"740A4661",X"6D696C79",X"3A205472",X"696F6E0A",X"44657669",X"63653A20",X"54384638",X"310A5769",X"6474683A",X"20310A50",X"41444445",
X"445F4249",X"54533A20",X"300A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",
X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",
X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"0A0A0A0A",X"168A2236",X"FFFE0740",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00010000",X"00000001",
X"00000000",X"00000000",X"00358341",X"50100060",X"00152200",X"002AC855",X"90AB2156",X"42AC8559",X"08311564",X"2AC85590",X"AB215642",
X"AC85590A",X"B2106220",X"4C559083",X"1106220C",X"44188831",X"10622AC8",X"5590AB21",X"5642AC85",X"590AB215",X"642AC851",X"90813146",
X"429CB002",X"60E4F041",X"88A32156",X"420C4559",X"0AB21564",X"2AC85590",X"AB215642",X"AC84098A",X"B2156420",X"A0559082",X"81026206",
X"C40D8AB2",X"00000000",X"00000000",X"00000000",X"90088082",X"40A09048",X"04122800",X"82410090",X"48241201",X"048A4120",X"00090480",
X"41209049",X"64120904",X"82492090",X"48241209",X"04824122",X"00090482",X"41209020",X"24060904",X"82410090",X"08240605",X"01920922",
X"90090482",X"41021248",X"240A7114",X"88406290",X"48A41229",X"04924122",X"9009048A",X"41239049",X"14500824",X"96412080",X"48241209",
X"04020120",X"00090480",X"41229048",X"24120904",X"82412090",X"48044209",X"148A4B20",X"00090482",X"41209148",X"0C920904",X"82412090",
X"48240221",X"04824520",X"90090482",X"41209048",X"20120134",X"82112590",X"48041209",X"00824100",X"00000000",X"00000000",X"00000000",
X"00001000",X"00000000",X"10000102",X"00081000",X"00000002",X"00140000",X"00000000",X"80000000",X"80000000",X"00040000",X"00000000",
X"00000001",X"00000000",X"00000004",X"00000000",X"00002000",X"10000000",X"00081401",X"00000000",X"08140100",X"00006220",X"10000700",
X"00000050",X"001C0001",X"00000004",X"00070000",X"80820110",X"080A0008",X"00000000",X"00801005",X"00000010",X"80040000",X"00000000",
X"00000000",X"00088800",X"00100400",X"00000000",X"00000000",X"00400000",X"00000000",X"00000440",X"00000000",X"00000000",X"00000000",
X"04000210",X"00000000",X"00200000",X"01000010",X"00000000",X"00000000",X"00000000",X"90093490",X"49248209",X"24B2092C",X"92492592",
X"C9E41209",X"14824121",X"00092482",X"49259048",X"24120904",X"80412090",X"48241209",X"04824125",X"00090482",X"41209049",X"C4B23824",
X"12412190",X"49224249",X"34820B20",X"90090496",X"41020148",X"0C824824",X"82052612",X"48248229",X"00024124",X"90082482",X"49209018",
X"1450432C",X"15052092",X"C8241079",X"048A4F20",X"00432482",X"45109048",X"04520904",X"924AA290",X"48241209",X"00924120",X"0009044A",
X"41209028",X"A492092A",X"82412090",X"49441271",X"241E4920",X"90090482",X"41209248",X"2490A82C",X"824B0090",X"C8245209",X"041A4B26",
X"00000000",X"00000000",X"00000000",X"0000100A",X"04020540",X"80002000",X"08000001",X"00800000",X"00000002",X"00000000",X"04020000",
X"00000000",X"02000000",X"00000000",X"00000002",X"00000000",X"00000000",X"00402110",X"48000200",X"00000420",X"00004000",X"00000000",
X"00042000",X"00402110",X"00000281",X"00000000",X"04200002",X"00005000",X"04040000",X"00022000",X"08400000",X"00000220",X"00000000",
X"00501000",X"00000000",X"10000000",X"00000000",X"00000000",X"00080000",X"00000000",X"00000200",X"00400010",X"00000000",X"00A00022",
X"10480000",X"00000000",X"00000000",X"00400100",X"00002001",X"00000020",X"00080002",X"00000000",X"00000000",X"00000000",X"00008000",
X"00000000",X"00000008",X"00000100",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000100",X"08402000",X"00000200",X"00800000",X"10000000",X"00000004",X"000A0101",X"00040000",X"000C0000",X"00000400",
X"00020000",X"00000000",X"01090000",X"00804008",X"08000000",X"80000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000400",
X"00004040",X"01000400",X"00000000",X"00020100",X"00400010",X"08000000",X"00000020",X"40000000",X"00000000",X"00000000",X"00200000",
X"00000000",X"00000000",X"00000C00",X"00000000",X"00000000",X"00000000",X"00000000",X"00000100",X"00000000",X"00000000",X"00800000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00050200",X"00204000",X"14000400",
X"010000D0",X"48000000",X"00000000",X"000C0580",X"00800000",X"000C0200",X"00000000",X"20080000",X"00001000",X"00080200",X"00002000",
X"100C0000",X"0000A000",X"20000000",X"00000000",X"00000200",X"01000000",X"00000000",X"02012000",X"00080800",X"00000000",X"000D0480",
X"00A00028",X"34000000",X"00018050",X"40000000",X"00000000",X"00040200",X"00800000",X"10000000",X"00000000",X"00080200",X"00000000",
X"00000000",X"00000000",X"048CC86C",X"92190C92",X"41209068",X"64120D04",X"A2412094",X"48241209",X"00004824",X"32090482",X"41209048",
X"24120904",X"82412090",X"48241209",X"00004824",X"120944A3",X"41A890C8",X"64138904",X"A2512194",X"68643A09",X"04804834",X"12A95F83",
X"493594CD",X"25769924",X"82413090",X"48741219",X"0480C824",X"32090482",X"6B21906A",X"A59A0906",X"82412890",X"4E271A0D",X"00024825",
X"12890482",X"59209048",X"241A0904",X"90188090",X"4A251209",X"00004A24",X"12400242",X"43209049",X"24120904",X"80012800",X"5A241209",
X"04804824",X"12090482",X"432890C8",X"241A0904",X"82512090",X"4AE41389",X"00000000",X"00000000",X"00000000",X"0008C080",X"6022000C",
X"08C00200",X"88004000",X"00000008",X"10000000",X"00000000",X"40000000",X"00000000",X"00600000",X"00000000",X"00000000",X"00000000",
X"00000050",X"00902000",X"00000000",X"4000020A",X"60888000",X"00000100",X"00003610",X"06122814",X"02042018",X"00001000",X"00100020",
X"00000000",X"0008000C",X"24450380",X"00080020",X"00000000",X"0000804C",X"00018002",X"04000000",X"00000000",X"00803000",X"0269A460",
X"00C00000",X"00000000",X"000926C0",X"04000000",X"00000000",X"024010B1",X"90000000",X"00000000",X"00000000",X"02000230",X"00804000",
X"00200000",X"04088030",X"00000000",X"00000000",X"00000000",X"9001201C",X"0F209148",X"0172082C",X"00C40700",X"49845214",X"11814122",
X"0000008A",X"45008110",X"20625824",X"88C10820",X"48A41229",X"00164100",X"0004820A",X"41208500",X"89457100",X"8E042284",X"42240604",
X"081CC412",X"90091002",X"01029049",X"A4404912",X"080F2031",X"4880E401",X"10021122",X"9008101E",X"44229140",X"C048203A",X"000A2591",
X"4420A089",X"04000520",X"0002041E",X"01229008",X"94522911",X"94490290",X"49241200",X"04800F02",X"00025080",X"C4229110",X"01122404",
X"16212080",X"20219279",X"18084060",X"90090482",X"41208848",X"84420904",X"80152090",X"01404600",X"00281000",X"00000000",X"00000000",
X"00000000",X"00083850",X"4A000080",X"08C00100",X"40022000",X"00888021",X"00000004",X"00032C10",X"00100A88",X"01642010",X"040A0008",
X"00000050",X"00980010",X"00000040",X"00000242",X"40A04221",X"0C280001",X"00000000",X"90000084",X"00002180",X"4A110000",X"C0055020",
X"50480000",X"80D08252",X"09880004",X"0000A140",X"0C010209",X"E4E10908",X"20C00402",X"0101B050",X"20421000",X"00002898",X"40040011",
X"00A00028",X"00042400",X"00800003",X"0000AA10",X"00002900",X"08800208",X"00005080",X"20000010",X"01404000",X"31148000",X"00002800",
X"00000000",X"20100000",X"00880000",X"40A40004",X"21008510",X"00000000",X"00000000",X"00000000",X"90089282",X"11209048",X"04320284",
X"84000630",X"28245201",X"01824006",X"00030202",X"41209021",X"88A0050C",X"84004810",X"0964B259",X"04824205",X"00000402",X"41201009",
X"44A65810",X"824A0D02",X"0024A0E8",X"40964100",X"84003014",X"42093042",X"A2080900",X"984A4532",X"08240449",X"08324900",X"90010092",
X"4B250389",X"60D20069",X"4000A041",X"49101203",X"24824085",X"00003438",X"0B208349",X"92120902",X"824C2490",X"08041208",X"04840120",
X"00052C80",X"49161000",X"040A0829",X"82412090",X"0920A051",X"24124884",X"84002482",X"412092A9",X"24C64322",X"92486490",X"41500A41",
X"34148005",X"00000000",X"00000000",X"00000000",X"00002000",X"00000000",X"00400000",X"08210600",X"81000008",X"00080096",X"00000080",
X"00000005",X"84020018",X"08240080",X"10804020",X"00000480",X"00000020",X"00000220",X"904020A0",X"00040030",X"08004860",X"000C0410",
X"0000322A",X"05020000",X"00020004",X"10001001",X"00002080",X"11000C20",X"00040408",X"00001320",X"02C00810",X"0A000012",X"00010000",
X"1000000A",X"00049818",X"04001300",X"80000000",X"08008200",X"40200000",X"80082000",X"00000002",X"04068044",X"10000090",X"00000000",
X"20C09100",X"10840010",X"00088000",X"00000000",X"80402010",X"080C0200",X"00400020",X"188020A0",X"00000000",X"00000000",X"00000000",
X"0001C0E6",X"44201008",X"3F420540",X"8FE5A1DC",X"88C4420D",X"16C84420",X"000DC0C8",X"402110CC",X"261EADC8",X"82F0ABD1",X"88840201",
X"10E845B9",X"00075488",X"40203008",X"37320111",X"E841E3D5",X"FE8403A5",X"CBEC45A0",X"040304E3",X"75B91008",X"045B9106",X"EAE2B810",
X"18173301",X"04804422",X"000DD6A6",X"6038306E",X"A43BBDD4",X"8B71A810",X"08264381",X"008471BA",X"000DC888",X"D0221008",X"37020106",
X"E0402010",X"0804022D",X"C083E020",X"000DC088",X"4020106E",X"84622DC6",X"E3702011",X"6E554A83",X"06EC4538",X"040DC080",X"4020DC08",
X"04022100",X"80422011",X"4C664203",X"18C45031",X"00000000",X"00000000",X"00000000",X"028CC00A",X"0E000000",X"00200000",X"10238200",
X"01008000",X"08440800",X"000C0644",X"080002A7",X"40901CC0",X"02000102",X"81008000",X"30640802",X"0004741C",X"0A050060",X"B3D06020",
X"640B87C1",X"E6400190",X"80540800",X"0000147B",X"33980280",X"0099C014",X"46201500",X"0153E070",X"04000800",X"028C8E3F",X"3C180066",
X"611994CC",X"0F358D00",X"0033D980",X"0000308B",X"0000C014",X"04070000",X"23000006",X"00000000",X"0000006C",X"E8032000",X"00047810",
X"00000027",X"03804446",X"633A0002",X"66915980",X"16740B98",X"00044000",X"0000CC00",X"00004000",X"00000003",X"4480C00C",X"E2623098",
X"00000000",X"00000000",X"00000000",X"0480C06B",X"14000000",X"38000CC0",X"03A062C1",X"1000000C",X"C7400000",X"00020140",X"00000010",
X"2A1C8000",X"02B1D8E0",X"00000000",X"006801B8",X"000F4660",X"00002050",X"031D8001",X"6000CAC8",X"76000584",X"43680190",X"44830663",
X"31502000",X"00058003",X"23A49800",X"10131D00",X"06600000",X"048CC702",X"201A2010",X"00000CC5",X"02F1CA20",X"00221982",X"000331D8",
X"0008C000",X"D0000000",X"3B000006",X"60044000",X"10000004",X"C003B000",X"000CC000",X"80000066",X"334004C1",X"03000000",X"36150882",
X"02600158",X"448CC000",X"00000010",X"00000201",X"00004000",X"0C0C0402",X"02202158",X"00000000",X"00000000",X"00000000",X"000CD6E7",
X"10000000",X"300009A0",X"802998E2",X"000C2000",X"C0540E00",X"000C06C4",X"00241233",X"33102220",X"020910EF",X"00000001",X"08F043BD",
X"000E7518",X"00002035",X"9B803218",X"70408CC0",X"260001E2",X"20D00F74",X"00000578",X"00440209",X"443BD109",X"07201203",X"811FD820",
X"2D184221",X"000DC603",X"30182001",X"09C07CC6",X"63318C20",X"093719A0",X"0093BCCC",X"0002F082",X"AC250000",X"6B800006",X"00002000",
X"00008216",X"F0036C24",X"000C5004",X"06070215",X"BB800667",X"73880010",X"6F111DC1",X"0B780FDE",X"00056800",X"00000010",X"08003200",
X"10020010",X"C038C07F",X"F669BD1A",X"00000000",X"00000000",X"00000000",X"90009036",X"04229000",X"20048904",X"80004010",X"12640561",
X"0C880802",X"0008148A",X"40409288",X"88007200",X"8A4C8D93",X"08840621",X"10284000",X"00005480",X"80228804",X"A0423900",X"200B0C09",
X"2982E070",X"91002825",X"9100148A",X"15220900",X"01042910",X"8940062B",X"10247050",X"502214A0",X"9001149E",X"04220001",X"60C00801",
X"1A401213",X"00A04201",X"11084122",X"00046988",X"45002148",X"91A06900",X"96051090",X"48240508",X"30584024",X"00086488",X"0F240401",
X"41022424",X"81412601",X"081150E5",X"14801A0C",X"91080118",X"11208240",X"04F04114",X"10482620",X"40010049",X"28000427",X"00000000",
X"00000000",X"00000000",X"00082108",X"2A410010",X"04800000",X"001A1482",X"80800024",X"10001424",X"00002810",X"00050141",X"00042101",
X"10040002",X"91100012",X"24020100",X"00020000",X"40450021",X"00806004",X"014E0200",X"81D0C868",X"20010507",X"00006014",X"00048244",
X"20A24001",X"10000E01",X"0000C088",X"0A000005",X"00020008",X"00443048",X"82D20040",X"1C008403",X"03048000",X"08960004",X"00000006",
X"20A24001",X"10000E01",X"0000C088",X"0A000005",X"00020008",X"00443048",X"82D20040",X"1C008403",X"03048000",X"08960004",X"08960004",
X"20A24001",X"10000E01",X"0000C088",X"0A000005",X"00020008",X"00443048",X"82D20040",X"1C008403",X"03048000",X"08960004",X"08960004",
X"00100680",X"00C62001",X"10180000",X"00000001",X"1C0A0102",X"00003814",X"CC022048",X"00844040",X"00000104",X"10008020",X"08960004",X"08960004");
	  signal   USER_MEM              : RAM_MEM_2;
      signal   XI                    : X_REG;                                             -- This array is identical to XII and holds the GPRs
	  signal   XII                   : X_REG;                                             -- This array is identical to XI and holds the GPRs
	  signal   DATA_FORMAT           : DATA_F;                                            -- Integer format for loading
	  signal   DATA_FORMAT_2         : DATA_F;                                            -- Integer format for loading passed to Stage 4
      signal   PC                    : signed(31 downto 0)            := X"00000001";     -- PC Register
	  signal   ARG1                  : signed(31 downto 0)            := X"00000000";     -- Argument 1 for operation	  
      signal   ARG2                  : signed(31 downto 0)            := X"00000000";     -- Argument 2 for operation	
	  signal   ARG3                  : signed(31 downto 0)            := X"00000000";     -- Argument 3 for operation
	  signal   SHIFT_STEPS           : integer range 0 to 31          := 0;               -- Shift Steps	  
	  signal   INSTRUCTION           : std_logic_vector(31 downto 0)  := X"00000000";     -- Instruction holding Register
	  signal   DESTINATION           : std_logic_vector(4 downto 0)   := "00000";         -- Instruction holding Register
	  signal   GPR                   : std_logic_vector(4 downto 0)   := "00000";         -- General Purpose Register Index
	  signal   U_REG                 : std_logic_vector(31 downto 0)  := X"00000000";     -- Formated U Type Immediate Register
      signal   RES                   : signed(63 downto 0)            := to_signed(0,64); -- Result after the instruction execution
      signal   STAGE2_EN             : std_logic                      := '0';             -- Enable bit for Stage 2 in the Pipeline
      signal   STAGE3_EN             : std_logic                      := '0';             -- Enable bit for Stage 3 in the Pipeline
      signal   STAGE4_EN             : std_logic                      := '0';             -- Enable bit for Stage 4 in the Pipeline
	  signal   J_PP                  : std_logic                      := '0';             -- JALR post processing flag
	  signal   PC_WRITE              : std_logic                      := '0';             -- PC write flag for Stage 4
	  signal   MEM_STORE             : std_logic                      := '0';             -- Register or Memory store flag for Stage 4
	  signal   PC_WRITE_2            : std_logic                      := '0';             -- PC write flag for Stage 4
	  signal   REG_STORE_2           : std_logic                      := '0';             -- Register or Memory store flag for Stage 4
	  signal   LOAD_OP               : std_logic                      := '0';             -- Load instrunction flag for post-processing
	  signal   sys_RES               : std_logic                      := '0';             -- Sincronously asserted system Reset
	  signal   sinc_T1               : std_logic                      := '0';             -- Sinchronous Clock 1 
	  signal   sinc_T2               : std_logic                      := '0';             -- Sinchronous Clock 2 
	  signal   sinc_T3               : std_logic                      := '0';             -- Sinchronous Clock 3 
	  signal   LOAD_DATA             : signed(31 downto 0)            := to_signed(0,32); -- LOAD Data
	  signal   SAVE_ADDRESS          : signed(31 downto 0)            := to_signed(0,32); -- SAVE ADDRESS
	  signal   SAVE_DATA             : signed(31 downto 0)            := to_signed(0,32); -- SAVE DATA
--
      function SIGN_EXTENDED_I(a: in STD_LOGIC_VECTOR ) return STD_LOGIC_VECTOR is
        begin
	      if (a(31) = '1') then return( "111111111111111111111" & a(30 downto 20));
		  else return( "000000000000000000000" & a(30 downto 20));
		  end if;
        end function SIGN_EXTENDED_I;
-- 
      function SIGN_EXTENDED_J(a: in STD_LOGIC_VECTOR ) return STD_LOGIC_VECTOR is
        begin
	      if (a(31) = '1') then return( "1111111111111" & a(19 downto 12)& a(20)& a(30 downto 21));
		  else return( "0000000000000" & a(19 downto 12)& a(20)& a(30 downto 21));
		  end if;
        end function SIGN_EXTENDED_J;
--
      function SIGN_EXTENDED_S(a: in STD_LOGIC_VECTOR ) return STD_LOGIC_VECTOR is
        begin
	      if (a(31) = '1') then return( "111111111111111111111" & a(30 downto 25)&a(11 downto 7));
		  else return( "000000000000000000000" & a(30 downto 25)&a(11 downto 7));
		  end if;
        end function SIGN_EXTENDED_S;
--
      function SHIFTED_U(a: in STD_LOGIC_VECTOR ) return STD_LOGIC_VECTOR is
        begin
	      return(a(31 downto 12) & "000000000000");
        end function SHIFTED_U;
--
      function SIGN_EXTENDED_8(a: in SIGNED) return SIGNED is
        begin
	      if (a(7) = '1') then return("1111111111111111111111111" & a(6 downto 0));
		  else return("0000000000000000000000000" & a(6 downto 0));
		  end if;
        end function SIGN_EXTENDED_8;
--
      function SIGN_EXTENDED_16(a: in SIGNED ) return SIGNED is
        begin
	      if (a(15) = '1') then return("11111111111111111" & a(14 downto 0));
		  else return("00000000000000000" & a(14 downto 0));
		  end if;
        end function SIGN_EXTENDED_16;
--
      function ZERO_EXTENDED_8(a: in SIGNED ) return SIGNED is
        begin
		  return("000000000000000000000000" & a(7 downto 0));
        end function ZERO_EXTENDED_8;
--
      function ZERO_EXTENDED_16(a: in SIGNED ) return SIGNED is
        begin
		  return("0000000000000000" & a(15 downto 0));
        end function ZERO_EXTENDED_16;
--
      function SLT(a,b: in SIGNED ) return SIGNED is
        begin
		  if a < b then
		     return ("00000000000000000000000000000001");
		  else
		     return("00000000000000000000000000000000");
		  end if;
        end function SLT;
--
      function SLTU(a,b: in SIGNED ) return SIGNED is
        begin
		  if unsigned(a) < unsigned(b) then
		     return ("00000000000000000000000000000001");
		  else
		     return("00000000000000000000000000000000");
		  end if;
        end function SLTU;
--
    begin
--
-- Synchronously assertion and asynchronously de-assertion of the system Reset
SYNC_RES: process (CLK, RST)
begin
     if RST = '0' then
	    sys_RES <= '0';
		sinc_T1 <= '0';
		sinc_T2 <= '0';
		sinc_T3 <= '0';
     else -- RST = '1'
	    sinc_T1 <= '1';
		sinc_T2 <= sinc_T1;
		sinc_T3 <= sinc_T2;
		if sinc_T1 = '1' AND sinc_T2 = '1' AND sinc_T3 = '1' then
		    sys_RES <= '1';
		end if;
	 end if; -- RST
end process SYNC_RES;
--
--
--============================== PIPELINE STAGE 1 ===================================
--================================== FETCHING =======================================
--
Stage_1: process (CLK, sys_RES)
begin
--
  if sys_RES = '0' then
    INSTRUCTION <= X"00000000";
	PC <= X"00000001";
	STAGE2_EN <= '0';
  else -- sys_RES = '1'
		if rising_edge(CLK) then
            -- Reading the instruction
            INSTRUCTION <= PROG_MEM(to_integer(PC));
			-- Enables the Stage 2
		    STAGE2_EN <= '1';
			--
		    CONTR_OUT <= std_logic_vector(RES(31 downto 0));
--
		    if (PC_WRITE='0') then
			    PC <= PC + 1;                            -- Increases the Program Counter
		    else
			    PC <= RES(31 downto 1) & '0';            -- Ipdates the PC from Pipeline Stage 2
			end if;
--
		  end if; -- rising edge (CLK)
--
    end if; -- RST
--
end process Stage_1;
--
--
--
--============================== PIPELINE STAGE 2 ===================================
--================================== ENCODING =======================================
--
Stage_2: process (CLK, sys_RES, STAGE2_EN)
begin
--
  if sys_RES = '0' then
	STAGE3_EN <= '0';
	PC_WRITE <= '0';
  else -- sys_RES = '1'
		if rising_edge(CLK) and STAGE2_EN = '1' then
            -- Enables the Stage 3 at the very beginning of the programm (second instruction after Reset)			
		    STAGE3_EN <= '1';
			--
			DESTINATION <= INSTRUCTION(19 downto 15);
			-- writing to the Program Counter register is disabled, unless otherwise stated in any of the states below
			PC_WRITE <= '0'; 
			ARG1 <= XI(to_integer(unsigned(INSTRUCTION(19 downto 15))));
			ARG2 <= XII(to_integer(unsigned(INSTRUCTION(24 downto 20))));
			SHIFT_STEPS <= to_integer(XII(to_integer(unsigned(INSTRUCTION(24 downto 20))))(4 downto 0));
			OPERATION <= o_SUM;
		    case INSTRUCTION(6 downto 2) is  -- Encoding the operand
              when "00000"               =>  ---------------------------------------- LOAD opcode
			    ARG2 <= signed(sign_extended_I(INSTRUCTION));
				OPERATION <= o_LOAD;
			    case INSTRUCTION(14 downto 12) is -- Encoding func.3
				   when "000"            =>  ------------------------ LB
				                             DATA_FORMAT <= l_8;
				   when "001"            =>  ------------------------ LH
				                             DATA_FORMAT <= l_16;
				   when "010"            =>  ------------------------ LW
				                             DATA_FORMAT <= l_32;
				   when "100"            =>  ------------------------ LBU
				                             DATA_FORMAT <= l_8_U;
				   when "101"            =>  ------------------------ LHU
				                             DATA_FORMAT <= l_16_U;
				   when others           =>  NULL;
				end case;
              when "00011"               =>  --------------------------------------- MISC_MEM opcode
			    case INSTRUCTION(14 downto 12) is -- Encoding func.3
				   when "000"            =>  ------------------------ FENCE
				   when "001"            =>  ------------------------ FENCEI
				   when others           =>  NULL;
				end case;
			  when "00100"               =>  --------------------------------------- OP-IMM opcode
			    SHIFT_STEPS <= to_integer(unsigned(INSTRUCTION(24 downto 20)));
				ARG2 <= signed(sign_extended_I(INSTRUCTION));
			    case INSTRUCTION(14 downto 12) is -- Encoding func.3
				   when "000"            =>  ------------------------ ADDI
				                             OPERATION <= o_SUM;
				   when "001"            =>  ------------------------ SLLI
				                             OPERATION <= o_SHIFT_LEFT;
				   when "010"            =>  ------------------------ SLTI
				                             OPERATION <= o_SLT;
				   when "011"            =>  ------------------------ SLTIU
				                             OPERATION <= o_SLTU;
				   when "100"            =>  ------------------------ XORI
				                             OPERATION <= o_XOR;
				   when "101"            => 
				     case INSTRUCTION(30) is -- Encoding func.7
					   when '0'          =>  ------------------------ SRLI;
					                         OPERATION <= o_SHIFT_RIGHT;
					   when '1'          =>  ------------------------ SRAI;
					                         OPERATION <= o_SRA;
					   when others       =>  NULL;
					 end case;
				   when "110"            =>  ------------------------ ORI
				                             OPERATION <= o_OR;
				   when "111"            =>  ------------------------ ANDI
				                             OPERATION <= o_AND;
				   when others           =>  NULL;
				end case;
			  when "00101"               =>  ------------------------ AUIPC / OPCODE
											 ARG1 <= signed(shifted_U(INSTRUCTION));
											 ARG2 <= PC;
			  when "01000"               =>  --------------------------------------- STORE opcode
				OPERATION <= o_SAVE;
				ARG3 <= signed(sign_extended_S(INSTRUCTION));
			    case INSTRUCTION(14 downto 12) is
				   when "000"            =>  ------------------------ SB
				                             DATA_FORMAT <= l_8_U;
				   when "001"            =>  ------------------------ SH
				                             DATA_FORMAT <= l_16_U;
				   when "010"            =>  ------------------------ SW
				                             DATA_FORMAT <= l_32;
				   when others           =>  NULL;
				end case;
              when "01100"               =>  --------------------------------------- OP opcode
			          case INSTRUCTION(14 downto 12) is -- Encoding func.3
				         when "000"      => 
				           case INSTRUCTION(30) is -- Encoding func.7
					         when '0'    =>  ------------------------ ADD
							                 OPERATION <= o_SUM;
					         when '1'    =>  ------------------------ SUB
							                 OPERATION <= o_SUB;
					         when others =>  NULL;
					       end case;
				         when "001"      =>  ------------------------ SLL
						                     OPERATION <= o_SHIFT_LEFT;
				         when "010"      =>  ------------------------ SLT
						                     OPERATION <= o_SLT;
				         when "011"      =>  ------------------------ SLTU
						                     OPERATION <= o_SLTU;
				         when "100"      =>  ------------------------ XOR
						                     OPERATION <= o_XOR;
				         when "101"      => 
				           case INSTRUCTION(30) is -- Encoding func.7
					         when '0'    =>  ------------------------ SRL
							                 OPERATION <= o_SHIFT_RIGHT;
					         when '1'    =>  ------------------------ SRA
							                 OPERATION <= o_SRA;
					         when others =>  NULL;
					       end case;
				         when "110"      =>  ------------------------ OR
						                     OPERATION <= o_OR;
				         when "111"      =>  ------------------------ AND
						                     OPERATION <= o_AND;
				         when others     =>  NULL;
				      end case;
              when "01101"               =>  ------------------------ LUI / OPCODE
											 ARG1 <= signed(shifted_U(INSTRUCTION));
											 ARG2 <= (others => '0');
              when "11000"               =>  ---------------------------------------- BRANCH opcode
			    case INSTRUCTION(14 downto 12) is -- Encoding func.3
				   when "000"            =>  ------------------------ BEQ
				   when "001"            =>  ------------------------ BNE
				   when "100"            =>  ------------------------ BLT
				   when "101"            =>  ------------------------ BGE
				   when "110"            =>  ------------------------ BLTU
				   when "111"            =>  ------------------------ BGEU
				   when others           =>  NULL;
				end case;
              when "11001"               =>  ------------------------ JALR / OPCODE
											 ARG2 <= signed (sign_extended_I(INSTRUCTION));
              when "11011"               =>  ------------------------ JAL / OPCODE
											 ARG1 <= signed (sign_extended_J(INSTRUCTION));
                                             ARG2 <= PC;
			  when "11100"               =>  ---------------------------------------- SYSTEM opcode
			    case INSTRUCTION(14 downto 12) is -- Encoding func.3
				   when "000"            =>
				     case INSTRUCTION(25)is  -- Encoding func.7
					   when '0'          =>  ------------------------ ECALL
					   when '1'          =>  ------------------------ EBREAK
					   when others       =>  NULL;
					  end case;
				   when "001"            =>  ------------------------ CSRRW
				   when "010"            =>  ------------------------ CSRRS
				   when "011"            =>  ------------------------ CSRRC
				   when "101"            =>  ------------------------ CSRRWI
				   when "110"            =>  ------------------------ CSRRSI
				   when "111"            =>  ------------------------ CSRRCI
				   when others           =>  NULL;
				end case;
              when others                =>  NULL;
           end case;
            --
         end if; -- rising edge (CLK)
  end if; -- sys_RES
end process Stage_2;
--
--
--
--============================== PIPELINE STAGE 3 ===================================
--================================= EXECUTING =======================================
--
Stage_3: process (CLK, sys_RES, STAGE3_EN)
begin
--
  if sys_RES = '0' then
	STAGE4_EN <= '0';
  else  -- sys_RES = '1'
		 if rising_edge(CLK) and (STAGE3_EN='1') then
--
			-- Enables the Stage 4 of the pipeline
			STAGE4_EN <= '1'; 
			-- Passes the GPR index from Stage 2 to Stage 4
            GPR <= DESTINATION;
--
            MEM_STORE <= '0'; -- the instruction result is stored in a GPR by default
			LOAD_OP <= '0';   -- no Load Operation flag by default
			case OPERATION is
			  when o_SUM         => RES(31 downto 0) <= ARG1 + ARG2;
			  when o_SUB         => RES(31 downto 0) <= ARG1 - ARG2;
			  when o_SHIFT_LEFT  => RES(31 downto 0) <= shift_left(ARG1, SHIFT_STEPS);
			  when o_SHIFT_RIGHT => RES(31 downto 0) <= shift_right(ARG1, SHIFT_STEPS);
			  when o_SRA         => RES(31 downto 0) <= ARG1 sra SHIFT_STEPS;
			  when o_AND         => RES(31 downto 0) <= ARG1 and ARG2;
			  when o_OR          => RES(31 downto 0) <= ARG1 or ARG2;
			  when o_XOR         => RES(31 downto 0) <= ARG1 xor ARG2;
			  when o_SLT         => RES(31 downto 0) <= SLT(ARG1, ARG2);
			  when o_SLTU        => RES(31 downto 0) <= SLTU(ARG1, ARG2);
			  when o_LOAD        => LOAD_DATA <= signed(USER_MEM(to_integer(ARG1 + ARG2)));
                        			LOAD_OP <= '1';               -- sets the Load Operation flag for Stage 4
									DATA_FORMAT_2 <= DATA_FORMAT; -- Passes the Load format from Stage 2 to Stage 4
			  when o_SAVE        => MEM_STORE <= '1';             -- result is stored in the user RAM memory
			                        SAVE_ADDRESS <= ARG1 + ARG3;
									case DATA_FORMAT_2 is
			                           when l_32   =>  SAVE_DATA <= ARG2;
				                       when l_16_U =>  SAVE_DATA <= ZERO_EXTENDED_16(ARG2);
				                       when l_8_U  =>  SAVE_DATA <= ZERO_EXTENDED_8(ARG2);
				                       when others => NULL;
			                        end case;
			  when others        => NULL;
		    end case;
--
		  end if; -- rising edge (CLK)
--
  end if; -- sys_RES
--
end process Stage_3;
--
--
--                
--============================== PIPELINE STAGE 4 ===================================
--=================================== SAVING ========================================
Stage_4: process (CLK, sys_RES, STAGE4_EN)
begin
    if sys_RES = '1' then
		  if rising_edge(CLK) and STAGE4_EN = '1' then
		  --
            if (MEM_STORE = '0') then
			  if LOAD_OP = '0' then
			    XI(to_integer(unsigned(GPR))) <= RES(31 downto 0) when J_PP = '0' else RES(31 downto 1) & '0';
			    XII(to_integer(unsigned(GPR))) <= RES(31 downto 0) when J_PP = '0' else RES(31 downto 1) & '0';
			  else
			     case DATA_FORMAT_2 is
				   when l_32 =>
			           XI(to_integer(unsigned(GPR))) <= LOAD_DATA;
			           XII(to_integer(unsigned(GPR))) <= LOAD_DATA;
				   when l_16 =>
			           XI(to_integer(unsigned(GPR))) <= SIGN_EXTENDED_16(LOAD_DATA);
			           XII(to_integer(unsigned(GPR))) <= SIGN_EXTENDED_16(LOAD_DATA);
				   when l_8 =>
			           XI(to_integer(unsigned(GPR))) <= SIGN_EXTENDED_8(LOAD_DATA);
			           XII(to_integer(unsigned(GPR))) <= SIGN_EXTENDED_8(LOAD_DATA);
				   when l_16_U =>
			           XI(to_integer(unsigned(GPR))) <= ZERO_EXTENDED_16(LOAD_DATA);
			           XII(to_integer(unsigned(GPR))) <= ZERO_EXTENDED_16(LOAD_DATA);
				   when l_8_U =>
			           XI(to_integer(unsigned(GPR))) <= ZERO_EXTENDED_8(LOAD_DATA);
			           XII(to_integer(unsigned(GPR))) <= ZERO_EXTENDED_8(LOAD_DATA);
				   when others => NULL;
				 end case;
			  end if;
			else
			  USER_MEM(to_integer(unsigned(SAVE_ADDRESS))) <= std_logic_vector(SAVE_DATA);
            end if; -- REG_STORE
		  --
		  end if; -- rising edge (CLK)
    end if; -- sys_RES
end process Stage_4;
--
--
--
--
end Behavioral;
