
//
// Verific Verilog Description of module RISC_V_Core
//

module RISC_V_Core (RST, CLK, CONTR_OUT, PORT_A) /* verific EFX_ATTRIBUTE_NETLIST__TOP_IS_VHDL=TRUE */ ;
    input RST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    input CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    output [31:0]CONTR_OUT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    output [31:0]PORT_A /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    
    wire n500_2;
    wire n522_2;
    wire n523_2;
    wire n524_2;
    wire n521_2;
    wire n525_2;
    wire n574_2;
    wire n526_2;
    wire n541_2;
    wire n531_2;
    wire n520_2;
    wire n519_2;
    wire n518_2;
    wire n517_2;
    wire n516_2;
    wire n515_2;
    wire n514_2;
    wire n513_2;
    wire n1615_2;
    wire n1649_2;
    wire n540_2;
    wire n539_2;
    wire n538_2;
    wire n537_2;
    wire n530_2;
    wire n529_2;
    wire n528_2;
    wire n512_2;
    wire n511_2;
    wire n510_2;
    wire n509_2;
    wire n508_2;
    wire n507_2;
    wire n501_2;
    wire n502_2;
    wire n495_2;
    wire n503_2;
    wire n496_2;
    wire n543_2;
    wire n504_2;
    wire n544_2;
    wire n505_2;
    wire n545_2;
    wire n546_2;
    wire n547_2;
    wire n548_2;
    wire n549_2;
    wire n550_2;
    wire n551_2;
    wire n552_2;
    wire n553_2;
    wire n554_2;
    wire n555_2;
    wire n556_2;
    wire n557_2;
    wire n558_2;
    wire n559_2;
    wire n560_2;
    wire n561_2;
    wire n562_2;
    wire n563_2;
    wire n564_2;
    wire n565_2;
    wire n566_2;
    wire n567_2;
    wire n568_2;
    wire n569_2;
    wire n570_2;
    wire n571_2;
    wire n572_2;
    wire n573_2;
    wire n506_2;
    wire n497_2;
    wire n498_2;
    wire n499_2;
    wire n1603_2;
    wire n1602_2;
    wire n1601_2;
    wire n1600_2;
    wire n1599_2;
    wire n1598_2;
    wire n1597_2;
    wire n1596_2;
    wire n1595_2;
    wire n1594_2;
    wire n1593_2;
    wire n1592_2;
    wire n1591_2;
    wire n1590_2;
    wire n1589_2;
    wire n1588_2;
    wire n1587_2;
    wire n1586_2;
    wire n1585_2;
    wire n1584_2;
    wire n1574_2;
    
    wire \ARG2[26] , \ARG2[4] , \ARG2[3] , n8, n9, STAGE2_EN, \PC[0] , 
        STAGE3_EN, \ARG2[2] , \ARG2[5] , \ARG2[1] , \DESTINATION[0] , 
        \ARG1[0] , \ARG2[0] , \SHIFT_STEPS[0] , \OPERATION[0] , \DATA_FORMAT[0] , 
        \ARG3[0] , STAGE4_EN, \ARG2[6] , \ARG2[7] , \ARG2[8] , \ARG2[9] , 
        \ARG2[10] , \ARG2[11] , \ARG2[12] , n32, n33, \ARG2[13] , 
        \LOAD_DATA[4] , \LOAD_DATA[5] , \LOAD_DATA[6] , \LOAD_DATA[7] , 
        n39, n40, \ARG3[2] , \ARG3[3] , \ARG3[4] , \ARG3[5] , \ARG3[6] , 
        \ARG3[7] , \ARG3[8] , \ARG3[9] , \GPR[0] , MEM_STORE, LOAD_OP, 
        \SHIFT_STEPS[1] , \SHIFT_STEPS[2] , \SHIFT_STEPS[3] , \SHIFT_STEPS[4] , 
        \OPERATION[1] , \OPERATION[2] , \OPERATION[3] , \DATA_FORMAT[1] , 
        \DATA_FORMAT[2] , \ARG3[1] , \DATA_FORMAT_2[0] , \SAVE_ADDRESS[0] , 
        \SAVE_DATA[0] , \ARG2[14] , \ARG2[15] , n51834, n51830, \ARG2[16] , 
        \ARG2[17] , \ARG2[18] , \ARG2[19] , \ARG2[25] , \ARG2[24] , 
        \ARG2[31] , \ARG2[23] , \ARG2[30] , \PC[7] , \PC[11] , \PC[15] , 
        \PC[19] , \PC[23] , \PC[27] , \PC[31] , \PC[3] , \PC[6] , 
        \PC[10] , \PC[14] , \PC[18] , \PC[22] , \PC[26] , \PC[30] , 
        \ARG1[31] , \PC[2] , \ARG2[22] , \ARG1[30] , \PC[5] , \PC[9] , 
        \PC[13] , \PC[17] , \PC[21] , \PC[25] , \PC[29] , \ARG2[21] , 
        \ARG1[29] , \LOAD_DATA[0] , \LOAD_DATA[1] , \LOAD_DATA[2] , 
        \LOAD_DATA[3] , \PC[1] , \ARG1[28] , \PC[4] , \PC[8] , \PC[12] , 
        \PC[16] , \PC[20] , \PC[24] , \PC[28] , \ARG1[27] , \ARG1[26] , 
        \ARG1[25] , n51730, n51726, \ARG1[24] , \ARG1[23] , \ARG1[22] , 
        \ARG1[21] , \ARG1[20] , \ARG1[19] , \ARG1[18] , \ARG1[17] , 
        \ARG1[16] , \ARG1[15] , \ARG1[14] , \ARG1[13] , \ARG1[12] , 
        \ARG1[11] , \ARG1[10] , \ARG1[9] , \ARG1[8] , \ARG1[7] , \ARG1[6] , 
        \ARG1[5] , \ARG1[4] , \ARG1[3] , \ARG1[2] , \ARG1[1] , \DESTINATION[4] , 
        \DESTINATION[3] , \XII[0][0] , \DESTINATION[2] , \XII[1][0] , 
        \DESTINATION[1] , \XII[2][0] , \XII[3][0] , \XII[4][0] , \XII[5][0] , 
        \XII[6][0] , \XII[7][0] , \XII[8][0] , \XII[9][0] , \XII[10][0] , 
        \XII[11][0] , \XII[12][0] , \XII[13][0] , \XII[14][0] , \XII[15][0] , 
        \XII[16][0] , \XII[17][0] , \XII[18][0] , \XII[19][0] , \XII[20][0] , 
        \XII[21][0] , \XII[22][0] , \XII[23][0] , \XII[24][0] , \XII[25][0] , 
        \XII[26][0] , \XII[27][0] , \XII[28][0] , \XII[29][0] , \XII[30][0] , 
        \XII[31][0] , \ARG2[20] , \ARG2[29] , \ARG2[28] , \ARG2[27] , 
        n221, \RES[7]_2~FF_brt_20_brt_70_brt_133_q_pinv , \CutToMuxOpt_21/n7 , 
        \RES[4]_2~FF_brt_123_q_pinv , \RES[3]_2~FF_brt_120_q_pinv , \RES[18]_2~FF_brt_89_q_pinv , 
        \RES[20]_2~FF_brt_92_q_pinv , \RES[22]_2~FF_brt_41_brt_98_q_pinv , 
        \CutToMuxOpt_23/n7 , \RES[23]_2~FF_brt_45_brt_100_q_pinv , \RES[12]_2~FF_brt_78_brt_145_q_pinv , 
        \GPR[1] , \GPR[2] , \GPR[3] , \GPR[4] , \LOAD_DATA[12] , \LOAD_DATA[13] , 
        \LOAD_DATA[14] , \LOAD_DATA[15] , \LOAD_DATA[16] , \LOAD_DATA[17] , 
        \LOAD_DATA[18] , \LOAD_DATA[19] , \LOAD_DATA[20] , \LOAD_DATA[21] , 
        \LOAD_DATA[22] , \LOAD_DATA[23] , \LOAD_DATA[24] , \LOAD_DATA[25] , 
        \LOAD_DATA[26] , \LOAD_DATA[27] , \LOAD_DATA[28] , \LOAD_DATA[29] , 
        \LOAD_DATA[30] , \LOAD_DATA[31] , \DATA_FORMAT_2[1] , \DATA_FORMAT_2[2] , 
        \SAVE_ADDRESS[1] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[4] , 
        \SAVE_ADDRESS[5] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[8] , 
        \SAVE_ADDRESS[9] , \SAVE_DATA[1] , \SAVE_DATA[2] , \SAVE_DATA[3] , 
        \SAVE_DATA[4] , \SAVE_DATA[5] , \SAVE_DATA[6] , \SAVE_DATA[7] , 
        \SAVE_DATA[8] , \SAVE_DATA[9] , \SAVE_DATA[10] , \SAVE_DATA[11] , 
        \SAVE_DATA[12] , \SAVE_DATA[13] , \SAVE_DATA[14] , \SAVE_DATA[15] , 
        \SAVE_DATA[16] , \SAVE_DATA[17] , \SAVE_DATA[18] , \SAVE_DATA[19] , 
        \SAVE_DATA[20] , \SAVE_DATA[21] , \SAVE_DATA[22] , \SAVE_DATA[23] , 
        \SAVE_DATA[24] , \SAVE_DATA[25] , \SAVE_DATA[26] , \SAVE_DATA[27] , 
        \SAVE_DATA[28] , \SAVE_DATA[29] , \SAVE_DATA[30] , \SAVE_DATA[31] , 
        \XI[0][8] , \XI[0][9] , \XI[0][10] , \XI[0][11] , \XI[0][12] , 
        \XI[0][13] , \XI[0][14] , \XI[0][15] , \XI[0][16] , \XI[0][17] , 
        \XI[0][18] , \XI[0][19] , \XI[0][20] , \XI[0][21] , \XI[0][22] , 
        \XI[0][23] , \XI[0][24] , \XI[0][25] , \XI[0][26] , \XI[0][27] , 
        \XI[0][28] , \XI[0][29] , \XI[0][30] , \XI[0][31] , \XI[1][8] , 
        \XI[1][9] , \XI[1][10] , \XI[1][11] , \XI[1][12] , \XI[1][13] , 
        \XI[1][14] , \XI[1][15] , \XI[1][16] , \XI[1][17] , \XI[1][18] , 
        \XI[1][19] , \XI[1][20] , \XI[1][21] , \XI[1][22] , \XI[1][23] , 
        \XI[1][24] , \XI[1][25] , \XI[1][26] , \XI[1][27] , \XI[1][28] , 
        \XI[1][29] , \XI[1][30] , \XI[1][31] , \XI[2][8] , \XI[2][9] , 
        \XI[2][10] , \XI[2][11] , \XI[2][12] , \XI[2][13] , \XI[2][14] , 
        \XI[2][15] , \XI[2][16] , \XI[2][17] , \XI[2][18] , \XI[2][19] , 
        \XI[2][20] , \XI[2][21] , \XI[2][22] , \XI[2][23] , \XI[2][24] , 
        \XI[2][25] , \XI[2][26] , \XI[2][27] , \XI[2][28] , \XI[2][29] , 
        \XI[2][30] , \XI[2][31] , \XI[3][8] , \XI[3][9] , \XI[3][10] , 
        \XI[3][11] , \XI[3][12] , \XI[3][13] , \XI[3][14] , \XI[3][15] , 
        \XI[3][16] , \XI[3][17] , \XI[3][18] , \XI[3][19] , \XI[3][20] , 
        \XI[3][21] , \XI[3][22] , \XI[3][23] , \XI[3][24] , \XI[3][25] , 
        \XI[3][26] , \XI[3][27] , \XI[3][28] , \XI[3][29] , \XI[3][30] , 
        \XI[3][31] , \XI[4][8] , \XI[4][9] , \XI[4][10] , \XI[4][11] , 
        \XI[4][12] , \XI[4][13] , \XI[4][14] , \XI[4][15] , \XI[4][16] , 
        \XI[4][17] , \XI[4][18] , \XI[4][19] , \XI[4][20] , \XI[4][21] , 
        \XI[4][22] , \XI[4][23] , \XI[4][24] , \XI[4][25] , \XI[4][26] , 
        \XI[4][27] , \XI[4][28] , \XI[4][29] , \XI[4][30] , \XI[4][31] , 
        \XI[5][8] , \XI[5][9] , \XI[5][10] , \XI[5][11] , \XI[5][12] , 
        \XI[5][13] , \XI[5][14] , \XI[5][15] , \XI[5][16] , \XI[5][17] , 
        \XI[5][18] , \XI[5][19] , \XI[5][20] , \XI[5][21] , \XI[5][22] , 
        \XI[5][23] , \XI[5][24] , \XI[5][25] , \XI[5][26] , \XI[5][27] , 
        \XI[5][28] , \XI[5][29] , \XI[5][30] , \XI[5][31] , \XI[6][8] , 
        \XI[6][9] , \XI[6][10] , \XI[6][11] , \XI[6][12] , \XI[6][13] , 
        \XI[6][14] , \XI[6][15] , \XI[6][16] , \XI[6][17] , \XI[6][18] , 
        \XI[6][19] , \XI[6][20] , \XI[6][21] , \XI[6][22] , \XI[6][23] , 
        \XI[6][24] , \XI[6][25] , \XI[6][26] , \XI[6][27] , \XI[6][28] , 
        \XI[6][29] , \XI[6][30] , \XI[6][31] , \XI[7][8] , \XI[7][9] , 
        \XI[7][10] , \XI[7][11] , \XI[7][12] , \XI[7][13] , \XI[7][14] , 
        \XI[7][15] , \XI[7][16] , \XI[7][17] , \XI[7][18] , \XI[7][19] , 
        \XI[7][20] , \XI[7][21] , \XI[7][22] , \XI[7][23] , \XI[7][24] , 
        \XI[7][25] , \XI[7][26] , \XI[7][27] , \XI[7][28] , \XI[7][29] , 
        \XI[7][30] , \XI[7][31] , \XI[8][8] , \XI[8][9] , \XI[8][10] , 
        \XI[8][11] , \XI[8][12] , \XI[8][13] , \XI[8][14] , \XI[8][15] , 
        \XI[8][16] , \XI[8][17] , \XI[8][18] , \XI[8][19] , \XI[8][20] , 
        \XI[8][21] , \XI[8][22] , \XI[8][23] , \XI[8][24] , \XI[8][25] , 
        \XI[8][26] , \XI[8][27] , \XI[8][28] , \XI[8][29] , \XI[8][30] , 
        \XI[8][31] , \XI[9][8] , \XI[9][9] , \XI[9][10] , \XI[9][11] , 
        \XI[9][12] , \XI[9][13] , \XI[9][14] , \XI[9][15] , \XI[9][16] , 
        \XI[9][17] , \XI[9][18] , \XI[9][19] , \XI[9][20] , \XI[9][21] , 
        \XI[9][22] , \XI[9][23] , \XI[9][24] , \XI[9][25] , \XI[9][26] , 
        \XI[9][27] , \XI[9][28] , \XI[9][29] , \XI[9][30] , \XI[9][31] , 
        \XI[10][8] , \XI[10][9] , \XI[10][10] , \XI[10][11] , \XI[10][12] , 
        \XI[10][13] , \XI[10][14] , \XI[10][15] , \XI[10][16] , \XI[10][17] , 
        \XI[10][18] , \XI[10][19] , \XI[10][20] , \XI[10][21] , \XI[10][22] , 
        \XI[10][23] , \XI[10][24] , \XI[10][25] , \XI[10][26] , \XI[10][27] , 
        \XI[10][28] , \XI[10][29] , \XI[10][30] , \XI[10][31] , \XI[11][8] , 
        \XI[11][9] , \XI[11][10] , \XI[11][11] , \XI[11][12] , \XI[11][13] , 
        \XI[11][14] , \XI[11][15] , \XI[11][16] , \XI[11][17] , \XI[11][18] , 
        \XI[11][19] , \XI[11][20] , \XI[11][21] , \XI[11][22] , \XI[11][23] , 
        \XI[11][24] , \XI[11][25] , \XI[11][26] , \XI[11][27] , \XI[11][28] , 
        \XI[11][29] , \XI[11][30] , \XI[11][31] , \XI[12][8] , \XI[12][9] , 
        \XI[12][10] , \XI[12][11] , \XI[12][12] , \XI[12][13] , \XI[12][14] , 
        \XI[12][15] , \XI[12][16] , \XI[12][17] , \XI[12][18] , \XI[12][19] , 
        \XI[12][20] , \XI[12][21] , \XI[12][22] , \XI[12][23] , \XI[12][24] , 
        \XI[12][25] , \XI[12][26] , \XI[12][27] , \XI[12][28] , \XI[12][29] , 
        \XI[12][30] , \XI[12][31] , \XI[13][8] , \XI[13][9] , \XI[13][10] , 
        \XI[13][11] , \XI[13][12] , \XI[13][13] , \XI[13][14] , \XI[13][15] , 
        \XI[13][16] , \XI[13][17] , \XI[13][18] , \XI[13][19] , \XI[13][20] , 
        \XI[13][21] , \XI[13][22] , \XI[13][23] , \XI[13][24] , \XI[13][25] , 
        \XI[13][26] , \XI[13][27] , \XI[13][28] , \XI[13][29] , \XI[13][30] , 
        \XI[13][31] , \XI[14][8] , \XI[14][9] , \XI[14][10] , \XI[14][11] , 
        \XI[14][12] , \XI[14][13] , \XI[14][14] , \XI[14][15] , \XI[14][16] , 
        \XI[14][17] , \XI[14][18] , \XI[14][19] , \XI[14][20] , \XI[14][21] , 
        \XI[14][22] , \XI[14][23] , \XI[14][24] , \XI[14][25] , \XI[14][26] , 
        \XI[14][27] , \XI[14][28] , \XI[14][29] , \XI[14][30] , \XI[14][31] , 
        \XI[15][8] , \XI[15][9] , \XI[15][10] , \XI[15][11] , \XI[15][12] , 
        \XI[15][13] , \XI[15][14] , \XI[15][15] , \XI[15][16] , \XI[15][17] , 
        \XI[15][18] , \XI[15][19] , \XI[15][20] , \XI[15][21] , \XI[15][22] , 
        \XI[15][23] , \XI[15][24] , \XI[15][25] , \XI[15][26] , \XI[15][27] , 
        \XI[15][28] , \XI[15][29] , \XI[15][30] , \XI[15][31] , \XI[16][8] , 
        \XI[16][9] , \XI[16][10] , \XI[16][11] , \XI[16][12] , \XI[16][13] , 
        \XI[16][14] , \XI[16][15] , \XI[16][16] , \XI[16][17] , \XI[16][18] , 
        \XI[16][19] , \XI[16][20] , \XI[16][21] , \XI[16][22] , \XI[16][23] , 
        \XI[16][24] , \XI[16][25] , \XI[16][26] , \XI[16][27] , \XI[16][28] , 
        \XI[16][29] , \XI[16][30] , \XI[16][31] , \XI[17][8] , \XI[17][9] , 
        \XI[17][10] , \XI[17][11] , \XI[17][12] , \XI[17][13] , \XI[17][14] , 
        \XI[17][15] , \XI[17][16] , \XI[17][17] , \XI[17][18] , \XI[17][19] , 
        \XI[17][20] , \XI[17][21] , \XI[17][22] , \XI[17][23] , \XI[17][24] , 
        \XI[17][25] , \XI[17][26] , \XI[17][27] , \XI[17][28] , \XI[17][29] , 
        \XI[17][30] , \XI[17][31] , \XI[18][8] , \XI[18][9] , \XI[18][10] , 
        \XI[18][11] , \XI[18][12] , \XI[18][13] , \XI[18][14] , \XI[18][15] , 
        \XI[18][16] , \XI[18][17] , \XI[18][18] , \XI[18][19] , \XI[18][20] , 
        \XI[18][21] , \XI[18][22] , \XI[18][23] , \XI[18][24] , \XI[18][25] , 
        \XI[18][26] , \XI[18][27] , \XI[18][28] , \XI[18][29] , \XI[18][30] , 
        \XI[18][31] , \XI[19][8] , \XI[19][9] , \XI[19][10] , \XI[19][11] , 
        \XI[19][12] , \XI[19][13] , \XI[19][14] , \XI[19][15] , \XI[19][16] , 
        \XI[19][17] , \XI[19][18] , \XI[19][19] , \XI[19][20] , \XI[19][21] , 
        \XI[19][22] , \XI[19][23] , \XI[19][24] , \XI[19][25] , \XI[19][26] , 
        \XI[19][27] , \XI[19][28] , \XI[19][29] , \XI[19][30] , \XI[19][31] , 
        \XI[20][8] , \XI[20][9] , \XI[20][10] , \XI[20][11] , \XI[20][12] , 
        \XI[20][13] , \XI[20][14] , \XI[20][15] , \XI[20][16] , \XI[20][17] , 
        \XI[20][18] , \XI[20][19] , \XI[20][20] , \XI[20][21] , \XI[20][22] , 
        \XI[20][23] , \XI[20][24] , \XI[20][25] , \XI[20][26] , \XI[20][27] , 
        \XI[20][28] , \XI[20][29] , \XI[20][30] , \XI[20][31] , \XI[21][8] , 
        \XI[21][9] , \XI[21][10] , \XI[21][11] , \XI[21][12] , \XI[21][13] , 
        \XI[21][14] , \XI[21][15] , \XI[21][16] , \XI[21][17] , \XI[21][18] , 
        \XI[21][19] , \XI[21][20] , \XI[21][21] , \XI[21][22] , \XI[21][23] , 
        \XI[21][24] , \XI[21][25] , \XI[21][26] , \XI[21][27] , \XI[21][28] , 
        \XI[21][29] , \XI[21][30] , \XI[21][31] , \XI[22][8] , \XI[22][9] , 
        \XI[22][10] , \XI[22][11] , \XI[22][12] , \XI[22][13] , \XI[22][14] , 
        \XI[22][15] , \XI[22][16] , \XI[22][17] , \XI[22][18] , \XI[22][19] , 
        \XI[22][20] , \XI[22][21] , \XI[22][22] , \XI[22][23] , \XI[22][24] , 
        \XI[22][25] , \XI[22][26] , \XI[22][27] , \XI[22][28] , \XI[22][29] , 
        \XI[22][30] , \XI[22][31] , \XI[23][8] , \XI[23][9] , \XI[23][10] , 
        \XI[23][11] , \XI[23][12] , \XI[23][13] , \XI[23][14] , \XI[23][15] , 
        \XI[23][16] , \XI[23][17] , \XI[23][18] , \XI[23][19] , \XI[23][20] , 
        \XI[23][21] , \XI[23][22] , \XI[23][23] , \XI[23][24] , \XI[23][25] , 
        \XI[23][26] , \XI[23][27] , \XI[23][28] , \XI[23][29] , \XI[23][30] , 
        \XI[23][31] , \XI[24][8] , \XI[24][9] , \XI[24][10] , \XI[24][11] , 
        \XI[24][12] , \XI[24][13] , \XI[24][14] , \XI[24][15] , \XI[24][16] , 
        \XI[24][17] , \XI[24][18] , \XI[24][19] , \XI[24][20] , \XI[24][21] , 
        \XI[24][22] , \XI[24][23] , \XI[24][24] , \XI[24][25] , \XI[24][26] , 
        \XI[24][27] , \XI[24][28] , \XI[24][29] , \XI[24][30] , \XI[24][31] , 
        \XI[25][8] , \XI[25][9] , \XI[25][10] , \XI[25][11] , \XI[25][12] , 
        \XI[25][13] , \XI[25][14] , \XI[25][15] , \XI[25][16] , \XI[25][17] , 
        \XI[25][18] , \XI[25][19] , \XI[25][20] , \XI[25][21] , \XI[25][22] , 
        \XI[25][23] , \XI[25][24] , \XI[25][25] , \XI[25][26] , \XI[25][27] , 
        \XI[25][28] , \XI[25][29] , \XI[25][30] , \XI[25][31] , \XI[26][8] , 
        \XI[26][9] , \XI[26][10] , \XI[26][11] , \XI[26][12] , \XI[26][13] , 
        \XI[26][14] , \XI[26][15] , \XI[26][16] , \XI[26][17] , \XI[26][18] , 
        \XI[26][19] , \XI[26][20] , \XI[26][21] , \XI[26][22] , \XI[26][23] , 
        \XI[26][24] , \XI[26][25] , \XI[26][26] , \XI[26][27] , \XI[26][28] , 
        \XI[26][29] , \XI[26][30] , \XI[26][31] , \XI[27][8] , \XI[27][9] , 
        \XI[27][10] , \XI[27][11] , \XI[27][12] , \XI[27][13] , \XI[27][14] , 
        \XI[27][15] , \XI[27][16] , \XI[27][17] , \XI[27][18] , \XI[27][19] , 
        \XI[27][20] , \XI[27][21] , \XI[27][22] , \XI[27][23] , \XI[27][24] , 
        \XI[27][25] , \XI[27][26] , \XI[27][27] , \XI[27][28] , \XI[27][29] , 
        \XI[27][30] , \XI[27][31] , \XI[28][8] , \XI[28][9] , \XI[28][10] , 
        \XI[28][11] , \XI[28][12] , \XI[28][13] , \XI[28][14] , \XI[28][15] , 
        \XI[28][16] , \XI[28][17] , \XI[28][18] , \XI[28][19] , \XI[28][20] , 
        \XI[28][21] , \XI[28][22] , \XI[28][23] , \XI[28][24] , \XI[28][25] , 
        \XI[28][26] , \XI[28][27] , \XI[28][28] , \XI[28][29] , \XI[28][30] , 
        \XI[28][31] , \XI[29][8] , \XI[29][9] , \XI[29][10] , \XI[29][11] , 
        \XI[29][12] , \XI[29][13] , \XI[29][14] , \XI[29][15] , \XI[29][16] , 
        \XI[29][17] , \XI[29][18] , \XI[29][19] , \XI[29][20] , \XI[29][21] , 
        \XI[29][22] , \XI[29][23] , \XI[29][24] , \XI[29][25] , \XI[29][26] , 
        \XI[29][27] , \XI[29][28] , \XI[29][29] , \XI[29][30] , \XI[29][31] , 
        \XI[30][8] , \XI[30][9] , \XI[30][10] , \XI[30][11] , \XI[30][12] , 
        \XI[30][13] , \XI[30][14] , \XI[30][15] , \XI[30][16] , \XI[30][17] , 
        \XI[30][18] , \XI[30][19] , \XI[30][20] , \XI[30][21] , \XI[30][22] , 
        \XI[30][23] , \XI[30][24] , \XI[30][25] , \XI[30][26] , \XI[30][27] , 
        \XI[30][28] , \XI[30][29] , \XI[30][30] , \XI[30][31] , \XI[31][8] , 
        \XI[31][9] , \XI[31][10] , \XI[31][11] , \XI[31][12] , \XI[31][13] , 
        \XI[31][14] , \XI[31][15] , \XI[31][16] , \XI[31][17] , \XI[31][18] , 
        \XI[31][19] , \XI[31][20] , \XI[31][21] , \XI[31][22] , \XI[31][23] , 
        \XI[31][24] , \XI[31][25] , \XI[31][26] , \XI[31][27] , \XI[31][28] , 
        \XI[31][29] , \XI[31][30] , \XI[31][31] , \XII[0][1] , \XII[0][2] , 
        \XII[0][3] , \XII[0][4] , \XII[0][5] , \XII[0][6] , \XII[0][7] , 
        \XII[1][1] , \XII[1][2] , \XII[1][3] , \XII[1][4] , \XII[1][5] , 
        \XII[1][6] , \XII[1][7] , \XII[2][1] , \XII[2][2] , \XII[2][3] , 
        \XII[2][4] , \XII[2][5] , \XII[2][6] , \XII[2][7] , \XII[3][1] , 
        \XII[3][2] , \XII[3][3] , \XII[3][4] , \XII[3][5] , \XII[3][6] , 
        \XII[3][7] , \XII[4][1] , \XII[4][2] , \XII[4][3] , \XII[4][4] , 
        \XII[4][5] , \XII[4][6] , \XII[4][7] , \XII[5][1] , \XII[5][2] , 
        \XII[5][3] , \XII[5][4] , \XII[5][5] , \XII[5][6] , \XII[5][7] , 
        \XII[6][1] , \XII[6][2] , \XII[6][3] , \XII[6][4] , \XII[6][5] , 
        \XII[6][6] , \XII[6][7] , \XII[7][1] , \XII[7][2] , \XII[7][3] , 
        \XII[7][4] , \XII[7][5] , \XII[7][6] , \XII[7][7] , \XII[8][1] , 
        \XII[8][2] , \XII[8][3] , \XII[8][4] , \XII[8][5] , \XII[8][6] , 
        \XII[8][7] , \XII[9][1] , \XII[9][2] , \XII[9][3] , \XII[9][4] , 
        \XII[9][5] , \XII[9][6] , \XII[9][7] , \XII[10][1] , \XII[10][2] , 
        \XII[10][3] , \XII[10][4] , \XII[10][5] , \XII[10][6] , \XII[10][7] , 
        \XII[11][1] , \XII[11][2] , \XII[11][3] , \XII[11][4] , \XII[11][5] , 
        \XII[11][6] , \XII[11][7] , \XII[12][1] , \XII[12][2] , \XII[12][3] , 
        \XII[12][4] , \XII[12][5] , \XII[12][6] , \XII[12][7] , \XII[13][1] , 
        \XII[13][2] , \XII[13][3] , \XII[13][4] , \XII[13][5] , \XII[13][6] , 
        \XII[13][7] , \XII[14][1] , \XII[14][2] , \XII[14][3] , \XII[14][4] , 
        \XII[14][5] , \XII[14][6] , \XII[14][7] , \XII[15][1] , \XII[15][2] , 
        \XII[15][3] , \XII[15][4] , \XII[15][5] , \XII[15][6] , \XII[15][7] , 
        \XII[16][1] , \XII[16][2] , \XII[16][3] , \XII[16][4] , \XII[16][5] , 
        \XII[16][6] , \XII[16][7] , \XII[17][1] , \XII[17][2] , \XII[17][3] , 
        \XII[17][4] , \XII[17][5] , \XII[17][6] , \XII[17][7] , \XII[18][1] , 
        \XII[18][2] , \XII[18][3] , \XII[18][4] , \XII[18][5] , \XII[18][6] , 
        \XII[18][7] , \XII[19][1] , \XII[19][2] , \XII[19][3] , \XII[19][4] , 
        \XII[19][5] , \XII[19][6] , \XII[19][7] , \XII[20][1] , \XII[20][2] , 
        \XII[20][3] , \XII[20][4] , \XII[20][5] , \XII[20][6] , \XII[20][7] , 
        \XII[21][1] , \XII[21][2] , \XII[21][3] , \XII[21][4] , \XII[21][5] , 
        \XII[21][6] , \XII[21][7] , \XII[22][1] , \XII[22][2] , \XII[22][3] , 
        \XII[22][4] , \XII[22][5] , \XII[22][6] , \XII[22][7] , \XII[23][1] , 
        \XII[23][2] , \XII[23][3] , \XII[23][4] , \XII[23][5] , \XII[23][6] , 
        \XII[23][7] , \XII[24][1] , \XII[24][2] , \XII[24][3] , \XII[24][4] , 
        \XII[24][5] , \XII[24][6] , \XII[24][7] , \XII[25][1] , \XII[25][2] , 
        \XII[25][3] , \XII[25][4] , \XII[25][5] , \XII[25][6] , \XII[25][7] , 
        \XII[26][1] , \XII[26][2] , \XII[26][3] , \XII[26][4] , \XII[26][5] , 
        \XII[26][6] , \XII[26][7] , \XII[27][1] , \XII[27][2] , \XII[27][3] , 
        \XII[27][4] , \XII[27][5] , \XII[27][6] , \XII[27][7] , \XII[28][1] , 
        \XII[28][2] , \XII[28][3] , \XII[28][4] , \XII[28][5] , \XII[28][6] , 
        \XII[28][7] , \XII[29][1] , \XII[29][2] , \XII[29][3] , \XII[29][4] , 
        \XII[29][5] , \XII[29][6] , \XII[29][7] , \XII[30][1] , \XII[30][2] , 
        \XII[30][3] , \XII[30][4] , \XII[30][5] , \XII[30][6] , \XII[30][7] , 
        \XII[31][1] , \XII[31][2] , \XII[31][3] , \XII[31][4] , \XII[31][5] , 
        \XII[31][6] , \XII[31][7] , n51738, n51734, \LOAD_DATA[8] , 
        \LOAD_DATA[9] , \LOAD_DATA[10] , \LOAD_DATA[11] , n51746, n51742, 
        n51754, n51750, n51762, n51758, n51770, n51766, n51778, 
        n51774, n51786, n51782, n51794, n51790, n51802, n51798, 
        n51810, n51806, n51818, n51814, n51826, n51822, n51842, 
        n51838, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
        n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
        n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
        n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, 
        n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
        n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
        n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
        n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, 
        n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
        n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
        n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
        n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
        n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
        n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
        n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
        n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
        n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
        n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, 
        n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, 
        n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
        n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
        n1508, n1509, n1510, n30664, \PC[0]__I , \INSTRUCTION[15] , 
        n49404, ceg_net35296, \INSTRUCTION[7] , n50065, n50476, n30807, 
        ceg_net408, \INSTRUCTION[9] , \INSTRUCTION[10] , \INSTRUCTION[11] , 
        \INSTRUCTION[25] , \INSTRUCTION[26] , \INSTRUCTION[27] , \INSTRUCTION[28] , 
        \INSTRUCTION[29] , n30678, n34248, n33468, n33460, ceg_net47657, 
        \INSTRUCTION[8] , n50605, ceg_net35302, \RES[2] , \CutToMuxOpt_19/n7 , 
        \RES[1] , \CutToMuxOpt_18/n7 , \CutToMuxOpt_22/n7 , \CutToMuxOpt_17/n7 , 
        \CutToMuxOpt_20/n7 , \RES[9]_2~FF_brt_0_q_pinv , \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_q_pinv , 
        \RES[15]_2~FF_brt_29_q_pinv , \CutToMuxOpt_16/n7 , \INSTRUCTION[19] , 
        \INSTRUCTION[18] , n19664, ceg_net27233, \INSTRUCTION[17] , 
        ceg_net27485, \INSTRUCTION[16] , ceg_net27737, ceg_net27989, 
        ceg_net28241, ceg_net28493, ceg_net28745, ceg_net28997, ceg_net29249, 
        ceg_net29501, ceg_net29753, ceg_net30005, ceg_net30257, ceg_net30509, 
        ceg_net30761, ceg_net31013, ceg_net31265, ceg_net31517, ceg_net31769, 
        ceg_net32021, ceg_net32273, ceg_net32525, ceg_net32777, ceg_net33029, 
        ceg_net33281, ceg_net33533, ceg_net33785, ceg_net34037, ceg_net34289, 
        ceg_net34541, ceg_net34793, ceg_net18979, \RES[13]_2~FF_brt_146_q_pinv , 
        n1795, n1614, n1613, n1612, n1611, n1610, n1609, n1608, 
        n1607, n1606, n1605, n1604, \RES[13]_2~FF_brt_147_q_pinv , 
        \RES[15]_2~FF_brt_30_brt_82_brt_151_q_pinv , \RES[19]_2~FF_brt_159_q_pinv , 
        \RES[22]_2~FF_brt_41_brt_97_brt_168_q_pinv , \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_q_pinv , 
        \RES[31]_2~FF_brt_66_brt_119_brt_191_q_pinv , \RES[0]_2~FF_brt_195_q , 
        \RES[0]_2~FF_brt_194_q , \RES[0]_2~FF_brt_193_q , \RES[0]_2~FF_brt_192_q , 
        \RES[31]_2~FF_brt_66_brt_119_brt_191_q , \RES[31]_2~FF_brt_66_brt_119_brt_190_q , 
        \RES[30]_2~FF_brt_189_q , \RES[30]_2~FF_brt_188_q , \RES[30]_2~FF_brt_187_q , 
        \RES[30]_2~FF_brt_186_q , \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185_q , 
        \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184_q , \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_q , 
        \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182_q , \RES[27]_2~FF_brt_55_brt_113_brt_181_q , 
        \RES[27]_2~FF_brt_55_brt_113_brt_180_q , \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179_q , 
        \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178_q , \RES[25]_2~FF_brt_108_brt_177_q , 
        \RES[25]_2~FF_brt_108_brt_176_q , \RES[25]_2~FF_brt_108_brt_175_q , 
        \RES[24]_2~FF_brt_49_brt_105_brt_174_q , \RES[24]_2~FF_brt_49_brt_105_brt_173_q , 
        \RES[24]_2~FF_brt_49_brt_105_brt_172_q , \RES[23]_2~FF_brt_45_brt_99_brt_171_q , 
        \RES[23]_2~FF_brt_45_brt_99_brt_170_q , \RES[22]_2~FF_brt_41_brt_97_brt_169_q , 
        \RES[22]_2~FF_brt_41_brt_97_brt_168_q , \RES[22]_2~FF_brt_41_brt_97_brt_167_q , 
        \RES[21]_2~FF_brt_96_brt_166_q , \RES[21]_2~FF_brt_96_brt_165_q , 
        \RES[20]_2~FF_brt_93_brt_164_q , \RES[20]_2~FF_brt_93_brt_163_q , 
        \RES[20]_2~FF_brt_93_brt_162_q , \RES[19]_2~FF_brt_161_q , \RES[19]_2~FF_brt_160_q , 
        n1575, n1573, n1572, n1571, n1570, n1569, n1568, n1567, 
        n1566, n1565, n1564, n1563, n1562, n1561, n1560, n1559, 
        n1558, n1557, n1556, n1555, n1554, n1553, n1552, n17577, 
        ceg_net41512, n17576, n17575, n17574, n17573, n17572, n17571, 
        n17570, n17569, ceg_net49709, n17568, n17567, n17566, n17565, 
        n17564, n17563, n17562, n17561, n17560, n17559, n17558, 
        n17557, n17556, n17555, n17554, n17610, ceg_net41704, n17609, 
        n17608, n17607, n17606, n17605, n17604, n17603, n17602, 
        ceg_net49773, n17601, n17600, n17599, n17598, n17597, n17596, 
        n17595, n17594, n17593, n17592, n17591, n17590, n17589, 
        n17588, n17587, n17643, ceg_net41896, n17642, n17641, n17640, 
        n17639, n17638, n17637, n17636, n17635, ceg_net49837, n17634, 
        n17633, n17632, n17631, n17630, n17629, n17628, n17627, 
        n17626, n17625, n17624, n17623, n17622, n17621, n17620, 
        n17676, ceg_net42088, n17675, n17674, n17673, n17672, n17671, 
        n17670, n17669, n17668, ceg_net49901, n17667, n17666, n17665, 
        n17664, n17663, n17662, n17661, n17660, n17659, n17658, 
        n17657, n17656, n17655, n17654, n17653, n17709, ceg_net42280, 
        n17708, n17707, n17706, n17705, n17704, n17703, n17702, 
        n17701, ceg_net49965, n17700, n17699, n17698, n17697, n17696, 
        n17695, n17694, n17693, n17692, n17691, n17690, n17689, 
        n17688, n17687, n17686, n17742, ceg_net42472, n17741, n17740, 
        n17739, n17738, n17737, n17736, n17735, n17734, ceg_net50029, 
        n17733, n17732, n17731, n17730, n17729, n17728, n17727, 
        n17726, n17725, n17724, n17723, n17722, n17721, n17720, 
        n17719, n17775, ceg_net42664, n17774, n17773, n17772, n17771, 
        n17770, n17769, n17768, n17767, ceg_net50093, n17766, n17765, 
        n17764, n17763, n17762, n17761, n17760, n17759, n17758, 
        n17757, n17756, n17755, n17754, n17753, n17752, n17808, 
        ceg_net42856, n17807, n17806, n17805, n17804, n17803, n17802, 
        n17801, n17800, ceg_net50157, n17799, n17798, n17797, n17796, 
        n17795, n17794, n17793, n17792, n17791, n17790, n17789, 
        n17788, n17787, n17786, n17785, n17841, ceg_net43048, n17840, 
        n17839, n17838, n17837, n17836, n17835, n17834, n17833, 
        ceg_net50221, n17832, n17831, n17830, n17829, n17828, n17827, 
        n17826, n17825, n17824, n17823, n17822, n17821, n17820, 
        n17819, n17818, n17874, ceg_net43240, n17873, n17872, n17871, 
        n17870, n17869, n17868, n17867, n17866, ceg_net50285, n17865, 
        n17864, n17863, n17862, n17861, n17860, n17859, n17858, 
        n17857, n17856, n17855, n17854, n17853, n17852, n17851, 
        n17907, ceg_net43432, n17906, n17905, n17904, n17903, n17902, 
        n17901, n17900, n17899, ceg_net50349, n17898, n17897, n17896, 
        n17895, n17894, n17893, n17892, n17891, n17890, n17889, 
        n17888, n17887, n17886, n17885, n17884, n17940, ceg_net43624, 
        n17939, n17938, n17937, n17936, n17935, n17934, n17933, 
        n17932, ceg_net50413, n17931, n17930, n17929, n17928, n17927, 
        n17926, n17925, n17924, n17923, n17922, n17921, n17920, 
        n17919, n17918, n17917, n17973, ceg_net43816, n17972, n17971, 
        n17970, n17969, n17968, n17967, n17966, n17965, ceg_net50477, 
        n17964, n17963, n17962, n17961, n17960, n17959, n17958, 
        n17957, n17956, n17955, n17954, n17953, n17952, n17951, 
        n17950, n18006, ceg_net44008, n18005, n18004, n18003, n18002, 
        n18001, n18000, n17999, n17998, ceg_net50541, n17997, n17996, 
        n17995, n17994, n17993, n17992, n17991, n17990, n17989, 
        n17988, n17987, n17986, n17985, n17984, n17983, n18039, 
        ceg_net44200, n18038, n18037, n18036, n18035, n18034, n18033, 
        n18032, n18031, ceg_net50605, n18030, n18029, n18028, n18027, 
        n18026, n18025, n18024, n18023, n18022, n18021, n18020, 
        n18019, n18018, n18017, n18016, n18072, ceg_net44392, n18071, 
        n18070, n18069, n18068, n18067, n18066, n18065, n18064, 
        ceg_net50669, n18063, n18062, n18061, n18060, n18059, n18058, 
        n18057, n18056, n18055, n18054, n18053, n18052, n18051, 
        n18050, n18049, n18105, ceg_net44584, n18104, n18103, n18102, 
        n18101, n18100, n18099, n18098, n18097, ceg_net50733, n18096, 
        n18095, n18094, n18093, n18092, n18091, n18090, n18089, 
        n18088, n18087, n18086, n18085, n18084, n18083, n18082, 
        n18138, ceg_net44776, n18137, n18136, n18135, n18134, n18133, 
        n18132, n18131, n18130, ceg_net50797, n18129, n18128, n18127, 
        n18126, n18125, n18124, n18123, n18122, n18121, n18120, 
        n18119, n18118, n18117, n18116, n18115, n18171, ceg_net44968, 
        n18170, n18169, n18168, n18167, n18166, n18165, n18164, 
        n18163, ceg_net50861, n18162, n18161, n18160, n18159, n18158, 
        n18157, n18156, n18155, n18154, n18153, n18152, n18151, 
        n18150, n18149, n18148, n18204, ceg_net45160, n18203, n18202, 
        n18201, n18200, n18199, n18198, n18197, n18196, ceg_net50925, 
        n18195, n18194, n18193, n18192, n18191, n18190, n18189, 
        n18188, n18187, n18186, n18185, n18184, n18183, n18182, 
        n18181, n18237, ceg_net45352, n18236, n18235, n18234, n18233, 
        n18232, n18231, n18230, n18229, ceg_net50989, n18228, n18227, 
        n18226, n18225, n18224, n18223, n18222, n18221, n18220, 
        n18219, n18218, n18217, n18216, n18215, n18214, n18270, 
        ceg_net45544, n18269, n18268, n18267, n18266, n18265, n18264, 
        n18263, n18262, ceg_net51053, n18261, n18260, n18259, n18258, 
        n18257, n18256, n18255, n18254, n18253, n18252, n18251, 
        n18250, n18249, n18248, n18247, n18303, ceg_net45736, n18302, 
        n18301, n18300, n18299, n18298, n18297, n18296, n18295, 
        ceg_net51117, n18294, n18293, n18292, n18291, n18290, n18289, 
        n18288, n18287, n18286, n18285, n18284, n18283, n18282, 
        n18281, n18280, n18336, ceg_net45928, n18335, n18334, n18333, 
        n18332, n18331, n18330, n18329, n18328, ceg_net51181, n18327, 
        n18326, n18325, n18324, n18323, n18322, n18321, n18320, 
        n18319, n18318, n18317, n18316, n18315, n18314, n18313, 
        n18369, ceg_net46120, n18368, n18367, n18366, n18365, n18364, 
        n18363, n18362, n18361, ceg_net51245, n18360, n18359, n18358, 
        n18357, n18356, n18355, n18354, n18353, n18352, n18351, 
        n18350, n18349, n18348, n18347, n18346, n18402, ceg_net46312, 
        n18401, n18400, n18399, n18398, n18397, n18396, n18395, 
        n18394, ceg_net51309, n18393, n18392, n18391, n18390, n18389, 
        n18388, n18387, n18386, n18385, n18384, n18383, n18382, 
        n18381, n18380, n18379, n18435, ceg_net46504, n18434, n18433, 
        n18432, n18431, n18430, n18429, n18428, n18427, ceg_net51373, 
        n18426, n18425, n18424, n18423, n18422, n18421, n18420, 
        n18419, n18418, n18417, n18416, n18415, n18414, n18413, 
        n18412, n18468, ceg_net46696, n18467, n18466, n18465, n18464, 
        n18463, n18462, n18461, n18460, ceg_net51437, n18459, n18458, 
        n18457, n18456, n18455, n18454, n18453, n18452, n18451, 
        n18450, n18449, n18448, n18447, n18446, n18445, n18501, 
        ceg_net46888, n18500, n18499, n18498, n18497, n18496, n18495, 
        n18494, n18493, ceg_net51501, n18492, n18491, n18490, n18489, 
        n18488, n18487, n18486, n18485, n18484, n18483, n18482, 
        n18481, n18480, n18479, n18478, n18534, ceg_net47080, n18533, 
        n18532, n18531, n18530, n18529, n18528, n18527, n18526, 
        ceg_net51565, n18525, n18524, n18523, n18522, n18521, n18520, 
        n18519, n18518, n18517, n18516, n18515, n18514, n18513, 
        n18512, n18511, n18567, ceg_net47272, n18566, n18565, n18564, 
        n18563, n18562, n18561, n18560, n18559, ceg_net51629, n18558, 
        n18557, n18556, n18555, n18554, n18553, n18552, n18551, 
        n18550, n18549, n18548, n18547, n18546, n18545, n18544, 
        n18600, ceg_net47464, n18599, n18598, n18597, n18596, n18595, 
        n18594, n18593, n18592, ceg_net51753, n18591, n18590, n18589, 
        n18588, n18587, n18586, n18585, n18584, n18583, n18582, 
        n18581, n18580, n18579, n18578, n18577, n19663, n19662, 
        n19661, n19660, n19659, n19658, n19657, \RES[19]_2~FF_brt_159_q , 
        \RES[18]_2~FF_brt_90_brt_157_q , \RES[18]_2~FF_brt_90_brt_156_q , 
        \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155_q , n2738, \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154_q , 
        n2741, \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153_q , \CutToMuxOpt_12/n7 , 
        n2744, \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152_q , n2747, \RES[15]_2~FF_brt_30_brt_82_brt_151_q , 
        n2750, \RES[14]_2~FF_brt_150_q , n2753, \RES[14]_2~FF_brt_149_q , 
        n2756, \RES[14]_2~FF_brt_148_q , n2759, \RES[13]_2~FF_brt_147_q , 
        n2762, \RES[13]_2~FF_brt_146_q , \CutToMuxOpt_11/n7 , n2765, 
        \RES[12]_2~FF_brt_78_brt_145_q , n2768, \RES[11]_2~FF_brt_144_q , 
        n2771, \RES[11]_2~FF_brt_143_q , n2774, \RES[11]_2~FF_brt_142_q , 
        n2777, \RES[11]_2~FF_brt_141_q , n2780, \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140_q , 
        n2783, \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139_q , \CutToMuxOpt_10/n7 , 
        n2786, \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q , n2789, \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q , 
        n2792, \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_q , n2795, \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135_q , 
        n2798, \RES[8]_2~FF_brt_21_brt_73_brt_134_q , n2801, \RES[7]_2~FF_brt_20_brt_70_brt_133_q , 
        n2804, \RES[7]_2~FF_brt_20_brt_70_brt_132_q , \CutToMuxOpt_9/n7 , 
        n2807, \RES[6]_2~FF_brt_131_q , n2810, \RES[6]_2~FF_brt_130_q , 
        n2813, \RES[6]_2~FF_brt_129_q , n2816, \RES[5]_2~FF_brt_128_q , 
        n2819, \RES[5]_2~FF_brt_127_q , n2822, \RES[5]_2~FF_brt_126_q , 
        n2825, \RES[4]_2~FF_brt_125_q , \CutToMuxOpt_8/n7 , \RES[4]_2~FF_brt_124_q , 
        \RES[4]_2~FF_brt_123_q , \RES[3]_2~FF_brt_121_q , \RES[3]_2~FF_brt_120_q , 
        \CutToMuxOpt_15/n7 , \RES[31]_2~FF_brt_66_brt_118_q , \RES[29]_2~FF_brt_16_brt_63_brt_116_q , 
        \RES[28]_2~FF_brt_15_brt_60_brt_114_q , \RES[27]_2~FF_brt_55_brt_112_q , 
        \RES[27]_2~FF_brt_55_brt_111_q , \RES[25]_2~FF_brt_109_q , \RES[25]_2~FF_brt_107_q , 
        \RES[25]_2~FF_brt_106_q , \RES[24]_2~FF_brt_49_brt_104_q , \RES[24]_2~FF_brt_49_brt_103_q , 
        \RES[24]_2~FF_brt_49_brt_102_q , \RES[23]_2~FF_brt_45_brt_100_q , 
        \CutToMuxOpt_14/n7 , \RES[22]_2~FF_brt_41_brt_98_q , \RES[21]_2~FF_brt_95_q , 
        \RES[21]_2~FF_brt_94_q , \CLK~O , \RES[20]_2~FF_brt_92_q , \RES[20]_2~FF_brt_91_q , 
        n5951, \RES[18]_2~FF_brt_89_q , \RES[18]_2~FF_brt_88_q , n5950, 
        \RES[17]_2~FF_brt_8_brt_37_brt_86_q , \RES[17]_2~FF_brt_8_brt_37_brt_85_q , 
        n5949, \RES[16]_2~FF_brt_5_brt_33_brt_83_q , n5948, \RES[15]_2~FF_brt_30_brt_81_q , 
        \RES[15]_2~FF_brt_30_brt_80_q , \RES[12]_2~FF_brt_79_q , n5947, 
        \RES[12]_2~FF_brt_77_q , n5946, \RES[10]_2~FF_brt_3_brt_28_brt_75_q , 
        n5945, n5944, \RES[8]_2~FF_brt_21_brt_72_q , \RES[8]_2~FF_brt_21_brt_71_q , 
        n5943, \RES[7]_2~FF_brt_20_brt_69_q , \RES[7]_2~FF_brt_20_brt_68_q , 
        \RES[31]_2~FF_brt_67_q , n5942, \RES[31]_2~FF_brt_65_q , \RES[31]_2~FF_brt_64_q , 
        n5941, \RES[29]_2~FF_brt_16_brt_62_q , \RES[29]_2~FF_brt_16_brt_61_q , 
        n5940, \RES[28]_2~FF_brt_15_brt_59_q , \RES[28]_2~FF_brt_15_brt_58_q , 
        \RES[28]_2~FF_brt_15_brt_57_q , \RES[27]_2~FF_brt_56_q , n5939, 
        \RES[27]_2~FF_brt_54_q , \RES[27]_2~FF_brt_53_q , n5938, \RES[26]_2~FF_brt_10_brt_51_q , 
        \RES[26]_2~FF_brt_10_brt_50_q , n5937, \RES[24]_2~FF_brt_48_q , 
        \RES[24]_2~FF_brt_47_q , \RES[24]_2~FF_brt_46_q , n5936, \RES[23]_2~FF_brt_44_q , 
        \RES[23]_2~FF_brt_43_q , \RES[23]_2~FF_brt_42_q , n5935, \CutToMuxOpt_13/n7 , 
        \RES[22]_2~FF_brt_39_q , \RES[22]_2~FF_brt_38_q , n5934, \RES[17]_2~FF_brt_8_brt_36_q , 
        \RES[17]_2~FF_brt_8_brt_35_q , \RES[17]_2~FF_brt_8_brt_34_q , n5933, 
        \RES[16]_2~FF_brt_5_brt_32_q , \RES[16]_2~FF_brt_5_brt_31_q , n5932, 
        \RES[15]_2~FF_brt_29_q , n5931, \RES[10]_2~FF_brt_3_brt_27_q , 
        n5930, \RES[9]_2~FF_brt_1_brt_25_q , \RES[9]_2~FF_brt_1_brt_24_q , 
        \RES[9]_2~FF_brt_1_brt_23_q , \RES[8]_2~FF_brt_22_q , n5929, n5928, 
        \RES[7]_2~FF_brt_19_q , \RES[7]_2~FF_brt_18_q , \RES[29]_2~FF_brt_17_q , 
        n5927, n5926, \RES[28]_2~FF_brt_14_q , \RES[28]_2~FF_brt_13_q , 
        \RES[26]_2~FF_brt_12_q , \RES[26]_2~FF_brt_11_q , n5925, \RES[17]_2~FF_brt_9_q , 
        n5924, \RES[17]_2~FF_brt_7_q , \RES[16]_2~FF_brt_6_q , n5923, 
        \RES[10]_2~FF_brt_4_q , n5922, n5921, \RES[9]_2~FF_brt_0_q , 
        n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, 
        n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
        n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
        n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, 
        n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
        n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
        n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3010, 
        n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
        n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
        n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
        n3037, n3038, n3041, n3042, n3043, n3044, n3045, n3046, 
        n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
        n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
        n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, 
        n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
        n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
        n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
        n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
        n3103, n3104, n3107, n3108, n3109, n3110, n3111, n3112, 
        n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, 
        n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
        n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
        n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, 
        n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
        n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, 
        n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, 
        n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
        n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
        n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
        n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, 
        n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
        n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
        n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, 
        n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, 
        n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
        n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, 
        n3251, n3252, n3255, n3256, n3257, n3258, n3259, n3260, 
        n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
        n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
        n3277, n3278, n3279, n3280, n3283, n3284, n3285, n3286, 
        n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
        n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
        n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, 
        n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, 
        n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
        n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
        n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
        n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, 
        n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
        n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, 
        n3371, n3372, n3375, n3376, n3377, n3378, n3379, n3380, 
        n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
        n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
        n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, 
        n3405, n3408, n3409, n3410, n3411, n3412, n3413, n3414, 
        n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
        n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, 
        n3431, n3432, n3433, n3434, n3435, n3438, n3439, n3440, 
        n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
        n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
        n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, 
        n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
        n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, 
        n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
        n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
        n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, 
        n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
        n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, 
        n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
        n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
        n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, 
        n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
        n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, 
        n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
        n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
        n3577, n3578, n3579, n3582, n3583, n3584, n3585, n3586, 
        n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, 
        n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
        n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3612, 
        n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, 
        n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, 
        n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, 
        n3637, n3638, n3639, n3642, n3643, n3644, n3645, n3646, 
        n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, 
        n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
        n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3672, 
        n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, 
        n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, 
        n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, 
        n3697, n3698, n3699, n3702, n3703, n3704, n3705, n3706, 
        n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, 
        n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
        n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3732, 
        n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, 
        n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, 
        n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, 
        n3757, n3758, n3759, n3762, n3763, n3764, n3765, n3766, 
        n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, 
        n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
        n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3792, 
        n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, 
        n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, 
        n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, 
        n3817, n3818, n3819, n3822, n3823, n3824, n3825, n3826, 
        n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, 
        n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
        n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3852, 
        n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, 
        n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, 
        n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, 
        n3877, n3878, n3879, n3882, n3883, n3884, n3885, n3886, 
        n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, 
        n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
        n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, 
        n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
        n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, 
        n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, 
        n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, 
        n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
        n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, 
        n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, 
        n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, 
        n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, 
        n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
        n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, 
        n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, 
        n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, 
        n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, 
        n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
        n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, 
        n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, 
        n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, 
        n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, 
        n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
        n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, 
        n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
        n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
        n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, 
        n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
        n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, 
        n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
        n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, 
        n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, 
        n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
        n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, 
        n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
        n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, 
        n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, 
        n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
        n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, 
        n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, 
        n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, 
        n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, 
        n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
        n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, 
        n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, 
        n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
        n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, 
        n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
        n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, 
        n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, 
        n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
        n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, 
        n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
        n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, 
        n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, 
        n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, 
        n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, 
        n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
        n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, 
        n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, 
        n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, 
        n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
        n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
        n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, 
        n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
        n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, 
        n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, 
        n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
        n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
        n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, 
        n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, 
        n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, 
        n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
        n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, 
        n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
        n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, 
        n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, 
        n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
        n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, 
        n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, 
        n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, 
        n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, 
        n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
        n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, 
        n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, 
        n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, 
        n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, 
        n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
        n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, 
        n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, 
        n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, 
        n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, 
        n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
        n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, 
        n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, 
        n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, 
        n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, 
        n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
        n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, 
        n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, 
        n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, 
        n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, 
        n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
        n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, 
        n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, 
        n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, 
        n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, 
        n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
        n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, 
        n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, 
        n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, 
        n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, 
        n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
        n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, 
        n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, 
        n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, 
        n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, 
        n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
        n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, 
        n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, 
        n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, 
        n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, 
        n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
        n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, 
        n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, 
        n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, 
        n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, 
        n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
        n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, 
        n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, 
        n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, 
        n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, 
        n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
        n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, 
        n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, 
        n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, 
        n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, 
        n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
        n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, 
        n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, 
        n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, 
        n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, 
        n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
        n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, 
        n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, 
        n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, 
        n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, 
        n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
        n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, 
        n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, 
        n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, 
        n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, 
        n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
        n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, 
        n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, 
        n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, 
        n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, 
        n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, 
        n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, 
        n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, 
        n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, 
        n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, 
        n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, 
        n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, 
        n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, 
        n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, 
        n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, 
        n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, 
        n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, 
        n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, 
        n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, 
        n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, 
        n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, 
        n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, 
        n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, 
        n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, 
        n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, 
        n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, 
        n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, 
        n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, 
        n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, 
        n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, 
        n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, 
        n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, 
        n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, 
        n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, 
        n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, 
        n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, 
        n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, 
        n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, 
        n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, 
        n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, 
        n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, 
        n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, 
        n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, 
        n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, 
        n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, 
        n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, 
        n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, 
        n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, 
        n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, 
        n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, 
        n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, 
        n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, 
        n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, 
        n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, 
        n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, 
        n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, 
        n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, 
        n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, 
        n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, 
        n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, 
        n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, 
        n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, 
        n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, 
        n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, 
        n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, 
        n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, 
        n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, 
        n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, 
        n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, 
        n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, 
        n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
        n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, 
        n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, 
        n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, 
        n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, 
        n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
        n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, 
        n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, 
        n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, 
        n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, 
        n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
        n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, 
        n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, 
        n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, 
        n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, 
        n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
        n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, 
        n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, 
        n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, 
        n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, 
        n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
        n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, 
        n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, 
        n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, 
        n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, 
        n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
        n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, 
        n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, 
        n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, 
        n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, 
        n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, 
        n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, 
        \CutToMuxOpt_7/n7 , \CutToMuxOpt_6/n7 , \CutToMuxOpt_5/n7 , \CutToMuxOpt_4/n7 , 
        \CutToMuxOpt_3/n7 , \CutToMuxOpt_2/n7 , \CutToMuxOpt_1/n7 , \CutToMuxOpt_0/n7 ;
    
    assign PORT_A[31] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[30] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[29] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[28] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[27] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[26] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[25] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[24] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[23] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[22] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[21] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[20] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[19] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[18] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[17] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[16] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[15] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[14] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[13] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[12] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[11] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[10] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[9] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[8] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE, EFX_ATTRIBUTE_PORT__IS_VHDL_PORT_NAME=TRUE */ ;
    assign PORT_A[0] = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 \CutToMuxOpt_11/Lut_0  (.I0(\XI[2][13] ), .I1(\XI[3][13] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_11/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_11/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_10/Lut_1  (.I0(\XI[0][12] ), .I1(\XI[1][12] ), 
            .I2(n2953), .I3(\CutToMuxOpt_10/n7 ), .O(n3408)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_10/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_10/Lut_0  (.I0(\XI[2][12] ), .I1(\XI[3][12] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_10/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_10/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_9/Lut_1  (.I0(\XI[0][11] ), .I1(\XI[1][11] ), 
            .I2(n2953), .I3(\CutToMuxOpt_9/n7 ), .O(n3375)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_9/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_9/Lut_0  (.I0(\XI[2][11] ), .I1(\XI[3][11] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_9/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_9/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_8/Lut_1  (.I0(\XI[0][10] ), .I1(\XI[1][10] ), 
            .I2(n2953), .I3(\CutToMuxOpt_8/n7 ), .O(n3339)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_8/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_8/Lut_0  (.I0(\XI[2][10] ), .I1(\XI[3][10] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_8/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_8/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_7/Lut_1  (.I0(\XI[0][9] ), .I1(\XI[1][9] ), .I2(n2953), 
            .I3(\CutToMuxOpt_7/n7 ), .O(n3313)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_7/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_7/Lut_0  (.I0(\XI[2][9] ), .I1(\XI[3][9] ), .I2(n2953), 
            .I3(n51770), .O(\CutToMuxOpt_7/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_7/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_6/Lut_1  (.I0(\XI[0][8] ), .I1(\XI[1][8] ), .I2(n2953), 
            .I3(\CutToMuxOpt_6/n7 ), .O(n3283)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_6/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_6/Lut_0  (.I0(\XI[2][8] ), .I1(\XI[3][8] ), .I2(n2953), 
            .I3(n51770), .O(\CutToMuxOpt_6/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_6/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_5/Lut_1  (.I0(\XII[0][7] ), .I1(\XII[1][7] ), 
            .I2(n2953), .I3(\CutToMuxOpt_5/n7 ), .O(n3255)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_5/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_5/Lut_0  (.I0(\XII[2][7] ), .I1(\XII[3][7] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_5/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_5/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_4/Lut_1  (.I0(\XII[0][6] ), .I1(\XII[1][6] ), 
            .I2(n2953), .I3(\CutToMuxOpt_4/n7 ), .O(n3227)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_4/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_4/Lut_0  (.I0(\XII[2][6] ), .I1(\XII[3][6] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_4/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_4/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \RES[4]_2~FF_brt_123_rtinv  (.I0(\RES[4]_2~FF_brt_123_q_pinv ), 
            .O(\RES[4]_2~FF_brt_123_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[4]_2~FF_brt_123_rtinv .LUTMASK = 16'h5555;
    EFX_FF \ARG2[26]~FF  (.D(n500_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[26]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[26]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[26]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[26]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[26]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[4]~FF  (.D(n522_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[4]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[4]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[4]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[4]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[4]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[3]~FF  (.D(n523_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[3]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[3]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[3]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[3]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[3]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[0]~FF  (.D(n1615_2), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[0]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[0]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[0]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[0]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[0]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[0]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \STAGE2_EN~FF  (.D(1'b1), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(STAGE2_EN)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \STAGE2_EN~FF .CLK_POLARITY = 1'b1;
    defparam \STAGE2_EN~FF .CE_POLARITY = 1'b1;
    defparam \STAGE2_EN~FF .SR_POLARITY = 1'b0;
    defparam \STAGE2_EN~FF .D_POLARITY = 1'b1;
    defparam \STAGE2_EN~FF .SR_SYNC = 1'b0;
    defparam \STAGE2_EN~FF .SR_VALUE = 1'b0;
    defparam \STAGE2_EN~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[0]~FF  (.D(\PC[0] ), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[0]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[0]~FF .CE_POLARITY = 1'b1;
    defparam \PC[0]~FF .SR_POLARITY = 1'b0;
    defparam \PC[0]~FF .D_POLARITY = 1'b0;
    defparam \PC[0]~FF .SR_SYNC = 1'b0;
    defparam \PC[0]~FF .SR_VALUE = 1'b0;
    defparam \PC[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \STAGE3_EN~FF  (.D(1'b1), .CE(STAGE2_EN), .CLK(\CLK~O ), .SR(n221), 
           .Q(STAGE3_EN)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \STAGE3_EN~FF .CLK_POLARITY = 1'b1;
    defparam \STAGE3_EN~FF .CE_POLARITY = 1'b1;
    defparam \STAGE3_EN~FF .SR_POLARITY = 1'b0;
    defparam \STAGE3_EN~FF .D_POLARITY = 1'b1;
    defparam \STAGE3_EN~FF .SR_SYNC = 1'b0;
    defparam \STAGE3_EN~FF .SR_VALUE = 1'b0;
    defparam \STAGE3_EN~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[2]~FF  (.D(n524_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[2]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[2]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[2]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[2]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[2]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[5]~FF  (.D(n521_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[5]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[5]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[5]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[5]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[5]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[1]~FF  (.D(n525_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[1]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[1]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[1]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[1]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[1]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DESTINATION[0]~FF  (.D(\INSTRUCTION[15] ), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DESTINATION[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DESTINATION[0]~FF .CLK_POLARITY = 1'b1;
    defparam \DESTINATION[0]~FF .CE_POLARITY = 1'b1;
    defparam \DESTINATION[0]~FF .SR_POLARITY = 1'b1;
    defparam \DESTINATION[0]~FF .D_POLARITY = 1'b1;
    defparam \DESTINATION[0]~FF .SR_SYNC = 1'b1;
    defparam \DESTINATION[0]~FF .SR_VALUE = 1'b0;
    defparam \DESTINATION[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[0]~FF  (.D(n574_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[0]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[0]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[0]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[0]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[0]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[0]~FF  (.D(n526_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[0]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[0]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[0]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[0]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[0]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SHIFT_STEPS[0]~FF  (.D(n541_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SHIFT_STEPS[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \SHIFT_STEPS[0]~FF .CLK_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[0]~FF .CE_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[0]~FF .SR_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[0]~FF .D_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[0]~FF .SR_SYNC = 1'b1;
    defparam \SHIFT_STEPS[0]~FF .SR_VALUE = 1'b0;
    defparam \SHIFT_STEPS[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \OPERATION[0]~FF  (.D(n531_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\OPERATION[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \OPERATION[0]~FF .CLK_POLARITY = 1'b1;
    defparam \OPERATION[0]~FF .CE_POLARITY = 1'b1;
    defparam \OPERATION[0]~FF .SR_POLARITY = 1'b1;
    defparam \OPERATION[0]~FF .D_POLARITY = 1'b1;
    defparam \OPERATION[0]~FF .SR_SYNC = 1'b1;
    defparam \OPERATION[0]~FF .SR_VALUE = 1'b0;
    defparam \OPERATION[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DATA_FORMAT[0]~FF  (.D(n49404), .CE(ceg_net35296), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DATA_FORMAT[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DATA_FORMAT[0]~FF .CLK_POLARITY = 1'b1;
    defparam \DATA_FORMAT[0]~FF .CE_POLARITY = 1'b0;
    defparam \DATA_FORMAT[0]~FF .SR_POLARITY = 1'b1;
    defparam \DATA_FORMAT[0]~FF .D_POLARITY = 1'b1;
    defparam \DATA_FORMAT[0]~FF .SR_SYNC = 1'b1;
    defparam \DATA_FORMAT[0]~FF .SR_VALUE = 1'b0;
    defparam \DATA_FORMAT[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[0]~FF  (.D(\INSTRUCTION[7] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[0]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[0]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[0]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[0]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[0]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[0]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \STAGE4_EN~FF  (.D(1'b1), .CE(STAGE3_EN), .CLK(\CLK~O ), .SR(n221), 
           .Q(STAGE4_EN)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \STAGE4_EN~FF .CLK_POLARITY = 1'b1;
    defparam \STAGE4_EN~FF .CE_POLARITY = 1'b1;
    defparam \STAGE4_EN~FF .SR_POLARITY = 1'b0;
    defparam \STAGE4_EN~FF .D_POLARITY = 1'b1;
    defparam \STAGE4_EN~FF .SR_SYNC = 1'b0;
    defparam \STAGE4_EN~FF .SR_VALUE = 1'b0;
    defparam \STAGE4_EN~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[6]~FF  (.D(n520_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[6]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[6]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[6]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[6]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[6]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[7]~FF  (.D(n519_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[7]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[7]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[7]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[7]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[7]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[8]~FF  (.D(n518_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[8]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[8]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[8]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[8]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[8]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[9]~FF  (.D(n517_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[9]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[9]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[9]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[9]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[9]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[10]~FF  (.D(n516_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[10]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[10]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[10]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[10]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[10]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[11]~FF  (.D(n515_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[11]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[11]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[11]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[11]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[11]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[12]~FF  (.D(n514_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[12]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[12]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[12]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[12]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[12]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[13]~FF  (.D(n513_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[13]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[13]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[13]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[13]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[13]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[9]_2~FF_brt_0_rtinv  (.I0(\RES[9]_2~FF_brt_0_q_pinv ), .O(\RES[9]_2~FF_brt_0_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[9]_2~FF_brt_0_rtinv .LUTMASK = 16'h5555;
    EFX_FF \ARG3[2]~FF  (.D(\INSTRUCTION[9] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[2]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[2]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[2]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[2]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[2]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[2]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[3]~FF  (.D(\INSTRUCTION[10] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[3]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[3]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[3]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[3]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[3]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[3]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[4]~FF  (.D(\INSTRUCTION[11] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[4]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[4]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[4]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[4]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[4]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[4]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[5]~FF  (.D(\INSTRUCTION[25] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[5]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[5]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[5]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[5]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[5]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[5]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[6]~FF  (.D(\INSTRUCTION[26] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[6]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[6]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[6]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[6]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[6]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[6]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[7]~FF  (.D(\INSTRUCTION[27] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[7]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[7]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[7]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[7]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[7]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[7]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[8]~FF  (.D(\INSTRUCTION[28] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[8]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[8]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[8]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[8]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[8]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[8]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[9]~FF  (.D(\INSTRUCTION[29] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[9]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[9]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[9]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[9]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[9]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[9]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \GPR[0]~FF  (.D(\DESTINATION[0] ), .CE(n30678), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\GPR[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \GPR[0]~FF .CLK_POLARITY = 1'b1;
    defparam \GPR[0]~FF .CE_POLARITY = 1'b1;
    defparam \GPR[0]~FF .SR_POLARITY = 1'b1;
    defparam \GPR[0]~FF .D_POLARITY = 1'b1;
    defparam \GPR[0]~FF .SR_SYNC = 1'b1;
    defparam \GPR[0]~FF .SR_VALUE = 1'b0;
    defparam \GPR[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MEM_STORE~FF  (.D(n34248), .CE(n30678), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(MEM_STORE)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \MEM_STORE~FF .CLK_POLARITY = 1'b1;
    defparam \MEM_STORE~FF .CE_POLARITY = 1'b1;
    defparam \MEM_STORE~FF .SR_POLARITY = 1'b1;
    defparam \MEM_STORE~FF .D_POLARITY = 1'b1;
    defparam \MEM_STORE~FF .SR_SYNC = 1'b1;
    defparam \MEM_STORE~FF .SR_VALUE = 1'b0;
    defparam \MEM_STORE~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LOAD_OP~FF  (.D(n1649_2), .CE(n30678), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(LOAD_OP)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \LOAD_OP~FF .CLK_POLARITY = 1'b1;
    defparam \LOAD_OP~FF .CE_POLARITY = 1'b1;
    defparam \LOAD_OP~FF .SR_POLARITY = 1'b1;
    defparam \LOAD_OP~FF .D_POLARITY = 1'b1;
    defparam \LOAD_OP~FF .SR_SYNC = 1'b1;
    defparam \LOAD_OP~FF .SR_VALUE = 1'b0;
    defparam \LOAD_OP~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SHIFT_STEPS[1]~FF  (.D(n540_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SHIFT_STEPS[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \SHIFT_STEPS[1]~FF .CLK_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[1]~FF .CE_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[1]~FF .SR_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[1]~FF .D_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[1]~FF .SR_SYNC = 1'b1;
    defparam \SHIFT_STEPS[1]~FF .SR_VALUE = 1'b0;
    defparam \SHIFT_STEPS[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SHIFT_STEPS[2]~FF  (.D(n539_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SHIFT_STEPS[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \SHIFT_STEPS[2]~FF .CLK_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[2]~FF .CE_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[2]~FF .SR_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[2]~FF .D_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[2]~FF .SR_SYNC = 1'b1;
    defparam \SHIFT_STEPS[2]~FF .SR_VALUE = 1'b0;
    defparam \SHIFT_STEPS[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SHIFT_STEPS[3]~FF  (.D(n538_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SHIFT_STEPS[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \SHIFT_STEPS[3]~FF .CLK_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[3]~FF .CE_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[3]~FF .SR_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[3]~FF .D_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[3]~FF .SR_SYNC = 1'b1;
    defparam \SHIFT_STEPS[3]~FF .SR_VALUE = 1'b0;
    defparam \SHIFT_STEPS[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SHIFT_STEPS[4]~FF  (.D(n537_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SHIFT_STEPS[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \SHIFT_STEPS[4]~FF .CLK_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[4]~FF .CE_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[4]~FF .SR_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[4]~FF .D_POLARITY = 1'b1;
    defparam \SHIFT_STEPS[4]~FF .SR_SYNC = 1'b1;
    defparam \SHIFT_STEPS[4]~FF .SR_VALUE = 1'b0;
    defparam \SHIFT_STEPS[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \OPERATION[1]~FF  (.D(n530_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\OPERATION[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \OPERATION[1]~FF .CLK_POLARITY = 1'b1;
    defparam \OPERATION[1]~FF .CE_POLARITY = 1'b1;
    defparam \OPERATION[1]~FF .SR_POLARITY = 1'b1;
    defparam \OPERATION[1]~FF .D_POLARITY = 1'b1;
    defparam \OPERATION[1]~FF .SR_SYNC = 1'b1;
    defparam \OPERATION[1]~FF .SR_VALUE = 1'b0;
    defparam \OPERATION[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \OPERATION[2]~FF  (.D(n529_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\OPERATION[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \OPERATION[2]~FF .CLK_POLARITY = 1'b1;
    defparam \OPERATION[2]~FF .CE_POLARITY = 1'b1;
    defparam \OPERATION[2]~FF .SR_POLARITY = 1'b1;
    defparam \OPERATION[2]~FF .D_POLARITY = 1'b1;
    defparam \OPERATION[2]~FF .SR_SYNC = 1'b1;
    defparam \OPERATION[2]~FF .SR_VALUE = 1'b0;
    defparam \OPERATION[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \OPERATION[3]~FF  (.D(n528_2), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\OPERATION[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \OPERATION[3]~FF .CLK_POLARITY = 1'b1;
    defparam \OPERATION[3]~FF .CE_POLARITY = 1'b1;
    defparam \OPERATION[3]~FF .SR_POLARITY = 1'b1;
    defparam \OPERATION[3]~FF .D_POLARITY = 1'b1;
    defparam \OPERATION[3]~FF .SR_SYNC = 1'b1;
    defparam \OPERATION[3]~FF .SR_VALUE = 1'b0;
    defparam \OPERATION[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DATA_FORMAT[1]~FF  (.D(n33468), .CE(ceg_net35296), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DATA_FORMAT[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DATA_FORMAT[1]~FF .CLK_POLARITY = 1'b1;
    defparam \DATA_FORMAT[1]~FF .CE_POLARITY = 1'b0;
    defparam \DATA_FORMAT[1]~FF .SR_POLARITY = 1'b1;
    defparam \DATA_FORMAT[1]~FF .D_POLARITY = 1'b1;
    defparam \DATA_FORMAT[1]~FF .SR_SYNC = 1'b1;
    defparam \DATA_FORMAT[1]~FF .SR_VALUE = 1'b0;
    defparam \DATA_FORMAT[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DATA_FORMAT[2]~FF  (.D(n33460), .CE(ceg_net47657), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DATA_FORMAT[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DATA_FORMAT[2]~FF .CLK_POLARITY = 1'b1;
    defparam \DATA_FORMAT[2]~FF .CE_POLARITY = 1'b0;
    defparam \DATA_FORMAT[2]~FF .SR_POLARITY = 1'b1;
    defparam \DATA_FORMAT[2]~FF .D_POLARITY = 1'b1;
    defparam \DATA_FORMAT[2]~FF .SR_SYNC = 1'b1;
    defparam \DATA_FORMAT[2]~FF .SR_VALUE = 1'b0;
    defparam \DATA_FORMAT[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG3[1]~FF  (.D(\INSTRUCTION[8] ), .CE(n50065), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\ARG3[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG3[1]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG3[1]~FF .CE_POLARITY = 1'b0;
    defparam \ARG3[1]~FF .SR_POLARITY = 1'b1;
    defparam \ARG3[1]~FF .D_POLARITY = 1'b1;
    defparam \ARG3[1]~FF .SR_SYNC = 1'b1;
    defparam \ARG3[1]~FF .SR_VALUE = 1'b0;
    defparam \ARG3[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DATA_FORMAT_2[0]~FF  (.D(\DATA_FORMAT[0] ), .CE(n50476), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DATA_FORMAT_2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \DATA_FORMAT_2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[0]~FF .CE_POLARITY = 1'b0;
    defparam \DATA_FORMAT_2[0]~FF .SR_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[0]~FF .D_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[0]~FF .SR_SYNC = 1'b1;
    defparam \DATA_FORMAT_2[0]~FF .SR_VALUE = 1'b0;
    defparam \DATA_FORMAT_2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[0]~FF  (.D(n32), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[0]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[0]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[0]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[0]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[0]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[0]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[0]~FF  (.D(\ARG2[0] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[0]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[0]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[0]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[0]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[0]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[14]~FF  (.D(n512_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[14]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[14]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[14]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[14]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[14]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[15]~FF  (.D(n511_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[15]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[15]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[15]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[15]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[15]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[16]~FF  (.D(n510_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[16]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[16]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[16]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[16]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[16]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[17]~FF  (.D(n509_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[17]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[17]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[17]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[17]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[17]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[18]~FF  (.D(n508_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[18]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[18]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[18]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[18]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[18]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[19]~FF  (.D(n507_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[19]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[19]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[19]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[19]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[19]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[25]~FF  (.D(n501_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[25]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[25]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[25]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[25]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[25]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[24]~FF  (.D(n502_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[24]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[24]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[24]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[24]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[24]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[31]~FF  (.D(n495_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[31]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[31]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[31]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[31]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[31]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[23]~FF  (.D(n503_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[23]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[23]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[23]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[23]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[23]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[30]~FF  (.D(n496_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[30]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[30]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[30]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[30]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[30]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[7]~FF  (.D(n1497), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[7]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[7]~FF .CE_POLARITY = 1'b1;
    defparam \PC[7]~FF .SR_POLARITY = 1'b0;
    defparam \PC[7]~FF .D_POLARITY = 1'b1;
    defparam \PC[7]~FF .SR_SYNC = 1'b0;
    defparam \PC[7]~FF .SR_VALUE = 1'b0;
    defparam \PC[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[11]~FF  (.D(n1489), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[11]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[11]~FF .CE_POLARITY = 1'b1;
    defparam \PC[11]~FF .SR_POLARITY = 1'b0;
    defparam \PC[11]~FF .D_POLARITY = 1'b1;
    defparam \PC[11]~FF .SR_SYNC = 1'b0;
    defparam \PC[11]~FF .SR_VALUE = 1'b0;
    defparam \PC[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[15]~FF  (.D(n1481), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[15]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[15]~FF .CE_POLARITY = 1'b1;
    defparam \PC[15]~FF .SR_POLARITY = 1'b0;
    defparam \PC[15]~FF .D_POLARITY = 1'b1;
    defparam \PC[15]~FF .SR_SYNC = 1'b0;
    defparam \PC[15]~FF .SR_VALUE = 1'b0;
    defparam \PC[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[19]~FF  (.D(n1473), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[19]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[19]~FF .CE_POLARITY = 1'b1;
    defparam \PC[19]~FF .SR_POLARITY = 1'b0;
    defparam \PC[19]~FF .D_POLARITY = 1'b1;
    defparam \PC[19]~FF .SR_SYNC = 1'b0;
    defparam \PC[19]~FF .SR_VALUE = 1'b0;
    defparam \PC[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[23]~FF  (.D(n1465), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[23]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[23]~FF .CE_POLARITY = 1'b1;
    defparam \PC[23]~FF .SR_POLARITY = 1'b0;
    defparam \PC[23]~FF .D_POLARITY = 1'b1;
    defparam \PC[23]~FF .SR_SYNC = 1'b0;
    defparam \PC[23]~FF .SR_VALUE = 1'b0;
    defparam \PC[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[27]~FF  (.D(n1457), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[27]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[27]~FF .CE_POLARITY = 1'b1;
    defparam \PC[27]~FF .SR_POLARITY = 1'b0;
    defparam \PC[27]~FF .D_POLARITY = 1'b1;
    defparam \PC[27]~FF .SR_SYNC = 1'b0;
    defparam \PC[27]~FF .SR_VALUE = 1'b0;
    defparam \PC[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[31]~FF  (.D(n1450), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[31]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[31]~FF .CE_POLARITY = 1'b1;
    defparam \PC[31]~FF .SR_POLARITY = 1'b0;
    defparam \PC[31]~FF .D_POLARITY = 1'b1;
    defparam \PC[31]~FF .SR_SYNC = 1'b0;
    defparam \PC[31]~FF .SR_VALUE = 1'b0;
    defparam \PC[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[2]~FF  (.D(\RES[2] ), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[2]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[2]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[2]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[2]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[2]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[2]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[6]~FF  (.D(n1609), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[6]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[6]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[6]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[6]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[6]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[6]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[10]~FF  (.D(n1605), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[10]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[10]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[10]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[10]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[10]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[10]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[14]~FF  (.D(n1601_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[14]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[14]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[14]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[14]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[14]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[14]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[18]~FF  (.D(n1597_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[18]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[18]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[18]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[18]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[18]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[18]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[22]~FF  (.D(n1593_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[22]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[22]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[22]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[22]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[22]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[22]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[26]~FF  (.D(n1589_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[26]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[26]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[26]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[26]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[26]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[26]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[30]~FF  (.D(n1585_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[30]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[30]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[30]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[30]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[30]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[30]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[3]~FF  (.D(n1505), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[3]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[3]~FF .CE_POLARITY = 1'b1;
    defparam \PC[3]~FF .SR_POLARITY = 1'b0;
    defparam \PC[3]~FF .D_POLARITY = 1'b1;
    defparam \PC[3]~FF .SR_SYNC = 1'b0;
    defparam \PC[3]~FF .SR_VALUE = 1'b0;
    defparam \PC[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[6]~FF  (.D(n1499), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[6]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[6]~FF .CE_POLARITY = 1'b1;
    defparam \PC[6]~FF .SR_POLARITY = 1'b0;
    defparam \PC[6]~FF .D_POLARITY = 1'b1;
    defparam \PC[6]~FF .SR_SYNC = 1'b0;
    defparam \PC[6]~FF .SR_VALUE = 1'b0;
    defparam \PC[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[10]~FF  (.D(n1491), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[10]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[10]~FF .CE_POLARITY = 1'b1;
    defparam \PC[10]~FF .SR_POLARITY = 1'b0;
    defparam \PC[10]~FF .D_POLARITY = 1'b1;
    defparam \PC[10]~FF .SR_SYNC = 1'b0;
    defparam \PC[10]~FF .SR_VALUE = 1'b0;
    defparam \PC[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[14]~FF  (.D(n1483), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[14]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[14]~FF .CE_POLARITY = 1'b1;
    defparam \PC[14]~FF .SR_POLARITY = 1'b0;
    defparam \PC[14]~FF .D_POLARITY = 1'b1;
    defparam \PC[14]~FF .SR_SYNC = 1'b0;
    defparam \PC[14]~FF .SR_VALUE = 1'b0;
    defparam \PC[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[18]~FF  (.D(n1475), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[18]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[18]~FF .CE_POLARITY = 1'b1;
    defparam \PC[18]~FF .SR_POLARITY = 1'b0;
    defparam \PC[18]~FF .D_POLARITY = 1'b1;
    defparam \PC[18]~FF .SR_SYNC = 1'b0;
    defparam \PC[18]~FF .SR_VALUE = 1'b0;
    defparam \PC[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[22]~FF  (.D(n1467), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[22]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[22]~FF .CE_POLARITY = 1'b1;
    defparam \PC[22]~FF .SR_POLARITY = 1'b0;
    defparam \PC[22]~FF .D_POLARITY = 1'b1;
    defparam \PC[22]~FF .SR_SYNC = 1'b0;
    defparam \PC[22]~FF .SR_VALUE = 1'b0;
    defparam \PC[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[26]~FF  (.D(n1459), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[26]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[26]~FF .CE_POLARITY = 1'b1;
    defparam \PC[26]~FF .SR_POLARITY = 1'b0;
    defparam \PC[26]~FF .D_POLARITY = 1'b1;
    defparam \PC[26]~FF .SR_SYNC = 1'b0;
    defparam \PC[26]~FF .SR_VALUE = 1'b0;
    defparam \PC[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[30]~FF  (.D(n1451), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[30]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[30]~FF .CE_POLARITY = 1'b1;
    defparam \PC[30]~FF .SR_POLARITY = 1'b0;
    defparam \PC[30]~FF .D_POLARITY = 1'b1;
    defparam \PC[30]~FF .SR_SYNC = 1'b0;
    defparam \PC[30]~FF .SR_VALUE = 1'b0;
    defparam \PC[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[31]~FF  (.D(n543_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[31]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[31]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[31]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[31]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[31]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[1]~FF  (.D(\RES[1] ), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[1]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[1]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[1]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[1]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[1]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[1]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[5]~FF  (.D(n1610), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[5]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[5]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[5]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[5]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[5]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[5]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[9]~FF  (.D(n1606), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[9]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[9]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[9]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[9]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[9]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[9]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[13]~FF  (.D(n1602_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[13]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[13]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[13]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[13]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[13]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[13]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[17]~FF  (.D(n1598_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[17]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[17]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[17]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[17]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[17]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[17]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[21]~FF  (.D(n1594_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[21]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[21]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[21]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[21]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[21]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[21]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[25]~FF  (.D(n1590_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[25]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[25]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[25]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[25]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[25]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[25]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[29]~FF  (.D(n1586_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[29]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[29]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[29]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[29]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[29]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[29]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[2]~FF  (.D(n1507), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[2]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[2]~FF .CE_POLARITY = 1'b1;
    defparam \PC[2]~FF .SR_POLARITY = 1'b0;
    defparam \PC[2]~FF .D_POLARITY = 1'b1;
    defparam \PC[2]~FF .SR_SYNC = 1'b0;
    defparam \PC[2]~FF .SR_VALUE = 1'b0;
    defparam \PC[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[22]~FF  (.D(n504_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[22]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[22]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[22]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[22]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[22]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[30]~FF  (.D(n544_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[30]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[30]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[30]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[30]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[30]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[5]~FF  (.D(n1501), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[5]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[5]~FF .CE_POLARITY = 1'b1;
    defparam \PC[5]~FF .SR_POLARITY = 1'b0;
    defparam \PC[5]~FF .D_POLARITY = 1'b1;
    defparam \PC[5]~FF .SR_SYNC = 1'b0;
    defparam \PC[5]~FF .SR_VALUE = 1'b0;
    defparam \PC[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[9]~FF  (.D(n1493), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[9]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[9]~FF .CE_POLARITY = 1'b1;
    defparam \PC[9]~FF .SR_POLARITY = 1'b0;
    defparam \PC[9]~FF .D_POLARITY = 1'b1;
    defparam \PC[9]~FF .SR_SYNC = 1'b0;
    defparam \PC[9]~FF .SR_VALUE = 1'b0;
    defparam \PC[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[13]~FF  (.D(n1485), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[13]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[13]~FF .CE_POLARITY = 1'b1;
    defparam \PC[13]~FF .SR_POLARITY = 1'b0;
    defparam \PC[13]~FF .D_POLARITY = 1'b1;
    defparam \PC[13]~FF .SR_SYNC = 1'b0;
    defparam \PC[13]~FF .SR_VALUE = 1'b0;
    defparam \PC[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[17]~FF  (.D(n1477), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[17]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[17]~FF .CE_POLARITY = 1'b1;
    defparam \PC[17]~FF .SR_POLARITY = 1'b0;
    defparam \PC[17]~FF .D_POLARITY = 1'b1;
    defparam \PC[17]~FF .SR_SYNC = 1'b0;
    defparam \PC[17]~FF .SR_VALUE = 1'b0;
    defparam \PC[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[21]~FF  (.D(n1469), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[21]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[21]~FF .CE_POLARITY = 1'b1;
    defparam \PC[21]~FF .SR_POLARITY = 1'b0;
    defparam \PC[21]~FF .D_POLARITY = 1'b1;
    defparam \PC[21]~FF .SR_SYNC = 1'b0;
    defparam \PC[21]~FF .SR_VALUE = 1'b0;
    defparam \PC[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[25]~FF  (.D(n1461), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[25]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[25]~FF .CE_POLARITY = 1'b1;
    defparam \PC[25]~FF .SR_POLARITY = 1'b0;
    defparam \PC[25]~FF .D_POLARITY = 1'b1;
    defparam \PC[25]~FF .SR_SYNC = 1'b0;
    defparam \PC[25]~FF .SR_VALUE = 1'b0;
    defparam \PC[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[29]~FF  (.D(n1453), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[29]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[29]~FF .CE_POLARITY = 1'b1;
    defparam \PC[29]~FF .SR_POLARITY = 1'b0;
    defparam \PC[29]~FF .D_POLARITY = 1'b1;
    defparam \PC[29]~FF .SR_SYNC = 1'b0;
    defparam \PC[29]~FF .SR_VALUE = 1'b0;
    defparam \PC[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[21]~FF  (.D(n505_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[21]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[21]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[21]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[21]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[21]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[29]~FF  (.D(n545_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[29]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[29]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[29]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[29]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[29]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[4]~FF  (.D(n1611), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[4]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[4]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[4]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[4]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[4]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[4]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[8]~FF  (.D(n1607), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[8]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[8]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[8]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[8]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[8]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[8]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[12]~FF  (.D(n1603_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[12]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[12]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[12]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[12]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[12]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[12]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[16]~FF  (.D(n1599_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[16]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[16]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[16]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[16]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[16]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[16]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[20]~FF  (.D(n1595_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[20]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[20]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[20]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[20]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[20]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[20]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[24]~FF  (.D(n1591_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[24]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[24]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[24]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[24]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[24]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[24]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[28]~FF  (.D(n1587_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[28]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[28]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[28]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[28]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[28]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[28]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[1]~FF  (.D(n1509), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[1]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[1]~FF .CE_POLARITY = 1'b1;
    defparam \PC[1]~FF .SR_POLARITY = 1'b0;
    defparam \PC[1]~FF .D_POLARITY = 1'b1;
    defparam \PC[1]~FF .SR_SYNC = 1'b0;
    defparam \PC[1]~FF .SR_VALUE = 1'b0;
    defparam \PC[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[28]~FF  (.D(n546_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[28]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[28]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[28]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[28]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[28]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[4]~FF  (.D(n1503), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[4]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[4]~FF .CE_POLARITY = 1'b1;
    defparam \PC[4]~FF .SR_POLARITY = 1'b0;
    defparam \PC[4]~FF .D_POLARITY = 1'b1;
    defparam \PC[4]~FF .SR_SYNC = 1'b0;
    defparam \PC[4]~FF .SR_VALUE = 1'b0;
    defparam \PC[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[8]~FF  (.D(n1495), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[8]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[8]~FF .CE_POLARITY = 1'b1;
    defparam \PC[8]~FF .SR_POLARITY = 1'b0;
    defparam \PC[8]~FF .D_POLARITY = 1'b1;
    defparam \PC[8]~FF .SR_SYNC = 1'b0;
    defparam \PC[8]~FF .SR_VALUE = 1'b0;
    defparam \PC[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[12]~FF  (.D(n1487), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[12]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[12]~FF .CE_POLARITY = 1'b1;
    defparam \PC[12]~FF .SR_POLARITY = 1'b0;
    defparam \PC[12]~FF .D_POLARITY = 1'b1;
    defparam \PC[12]~FF .SR_SYNC = 1'b0;
    defparam \PC[12]~FF .SR_VALUE = 1'b0;
    defparam \PC[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[16]~FF  (.D(n1479), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[16]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[16]~FF .CE_POLARITY = 1'b1;
    defparam \PC[16]~FF .SR_POLARITY = 1'b0;
    defparam \PC[16]~FF .D_POLARITY = 1'b1;
    defparam \PC[16]~FF .SR_SYNC = 1'b0;
    defparam \PC[16]~FF .SR_VALUE = 1'b0;
    defparam \PC[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[20]~FF  (.D(n1471), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[20]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[20]~FF .CE_POLARITY = 1'b1;
    defparam \PC[20]~FF .SR_POLARITY = 1'b0;
    defparam \PC[20]~FF .D_POLARITY = 1'b1;
    defparam \PC[20]~FF .SR_SYNC = 1'b0;
    defparam \PC[20]~FF .SR_VALUE = 1'b0;
    defparam \PC[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[24]~FF  (.D(n1463), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[24]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[24]~FF .CE_POLARITY = 1'b1;
    defparam \PC[24]~FF .SR_POLARITY = 1'b0;
    defparam \PC[24]~FF .D_POLARITY = 1'b1;
    defparam \PC[24]~FF .SR_SYNC = 1'b0;
    defparam \PC[24]~FF .SR_VALUE = 1'b0;
    defparam \PC[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PC[28]~FF  (.D(n1455), .CE(1'b1), .CLK(\CLK~O ), .SR(n221), 
           .Q(\PC[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \PC[28]~FF .CLK_POLARITY = 1'b1;
    defparam \PC[28]~FF .CE_POLARITY = 1'b1;
    defparam \PC[28]~FF .SR_POLARITY = 1'b0;
    defparam \PC[28]~FF .D_POLARITY = 1'b1;
    defparam \PC[28]~FF .SR_SYNC = 1'b0;
    defparam \PC[28]~FF .SR_VALUE = 1'b0;
    defparam \PC[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[27]~FF  (.D(n547_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[27]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[27]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[27]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[27]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[27]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[3]~FF  (.D(n1612), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[3]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[3]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[3]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[3]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[3]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[3]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[7]~FF  (.D(n1608), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[7]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[7]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[7]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[7]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[7]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[7]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[11]~FF  (.D(n1604), .CE(n221), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(CONTR_OUT[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[11]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[11]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[11]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[11]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[11]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[11]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[15]~FF  (.D(n1600_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[15]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[15]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[15]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[15]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[15]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[15]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[19]~FF  (.D(n1596_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[19]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[19]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[19]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[19]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[19]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[19]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[23]~FF  (.D(n1592_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[23]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[23]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[23]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[23]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[23]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[23]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[27]~FF  (.D(n1588_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[27]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[27]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[27]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[27]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[27]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[27]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CONTR_OUT[31]~FF  (.D(n1584_2), .CE(n221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(CONTR_OUT[31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(380)
    defparam \CONTR_OUT[31]~FF .CLK_POLARITY = 1'b1;
    defparam \CONTR_OUT[31]~FF .CE_POLARITY = 1'b1;
    defparam \CONTR_OUT[31]~FF .SR_POLARITY = 1'b1;
    defparam \CONTR_OUT[31]~FF .D_POLARITY = 1'b1;
    defparam \CONTR_OUT[31]~FF .SR_SYNC = 1'b1;
    defparam \CONTR_OUT[31]~FF .SR_VALUE = 1'b0;
    defparam \CONTR_OUT[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[26]~FF  (.D(n548_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[26]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[26]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[26]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[26]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[26]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[25]~FF  (.D(n549_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[25]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[25]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[25]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[25]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[25]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[24]~FF  (.D(n550_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[24]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[24]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[24]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[24]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[24]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[23]~FF  (.D(n551_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[23]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[23]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[23]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[23]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[23]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[22]~FF  (.D(n552_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[22]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[22]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[22]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[22]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[22]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[21]~FF  (.D(n553_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[21]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[21]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[21]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[21]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[21]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[20]~FF  (.D(n554_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[20]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[20]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[20]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[20]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[20]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[19]~FF  (.D(n555_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[19]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[19]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[19]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[19]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[19]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[18]~FF  (.D(n556_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[18]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[18]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[18]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[18]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[18]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[17]~FF  (.D(n557_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[17]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[17]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[17]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[17]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[17]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[16]~FF  (.D(n558_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[16]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[16]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[16]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[16]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[16]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[15]~FF  (.D(n559_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[15]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[15]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[15]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[15]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[15]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[14]~FF  (.D(n560_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[14]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[14]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[14]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[14]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[14]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[13]~FF  (.D(n561_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[13]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[13]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[13]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[13]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[13]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[12]~FF  (.D(n562_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[12]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[12]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[12]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[12]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[12]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[11]~FF  (.D(n563_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[11]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[11]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[11]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[11]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[11]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[10]~FF  (.D(n564_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[10]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[10]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[10]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[10]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[10]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[9]~FF  (.D(n565_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[9]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[9]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[9]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[9]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[9]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[8]~FF  (.D(n566_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[8]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[8]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[8]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[8]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[8]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[7]~FF  (.D(n567_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[7]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[7]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[7]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[7]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[7]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[6]~FF  (.D(n568_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[6]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[6]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[6]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[6]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[6]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[5]~FF  (.D(n569_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[5]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[5]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[5]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[5]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[5]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[4]~FF  (.D(n570_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[4]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[4]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[4]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[4]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[4]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[3]~FF  (.D(n571_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[3]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[3]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[3]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[3]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[3]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[2]~FF  (.D(n572_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[2]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[2]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[2]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[2]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[2]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG1[1]~FF  (.D(n573_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG1[1]~FF .CE_POLARITY = 1'b1;
    defparam \ARG1[1]~FF .SR_POLARITY = 1'b1;
    defparam \ARG1[1]~FF .D_POLARITY = 1'b1;
    defparam \ARG1[1]~FF .SR_SYNC = 1'b1;
    defparam \ARG1[1]~FF .SR_VALUE = 1'b0;
    defparam \ARG1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DESTINATION[4]~FF  (.D(\INSTRUCTION[19] ), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DESTINATION[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DESTINATION[4]~FF .CLK_POLARITY = 1'b1;
    defparam \DESTINATION[4]~FF .CE_POLARITY = 1'b1;
    defparam \DESTINATION[4]~FF .SR_POLARITY = 1'b1;
    defparam \DESTINATION[4]~FF .D_POLARITY = 1'b1;
    defparam \DESTINATION[4]~FF .SR_SYNC = 1'b1;
    defparam \DESTINATION[4]~FF .SR_VALUE = 1'b0;
    defparam \DESTINATION[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DESTINATION[3]~FF  (.D(\INSTRUCTION[18] ), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DESTINATION[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DESTINATION[3]~FF .CLK_POLARITY = 1'b1;
    defparam \DESTINATION[3]~FF .CE_POLARITY = 1'b1;
    defparam \DESTINATION[3]~FF .SR_POLARITY = 1'b1;
    defparam \DESTINATION[3]~FF .D_POLARITY = 1'b1;
    defparam \DESTINATION[3]~FF .SR_SYNC = 1'b1;
    defparam \DESTINATION[3]~FF .SR_VALUE = 1'b0;
    defparam \DESTINATION[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][0]~FF  (.D(n19664), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DESTINATION[2]~FF  (.D(\INSTRUCTION[17] ), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DESTINATION[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DESTINATION[2]~FF .CLK_POLARITY = 1'b1;
    defparam \DESTINATION[2]~FF .CE_POLARITY = 1'b1;
    defparam \DESTINATION[2]~FF .SR_POLARITY = 1'b1;
    defparam \DESTINATION[2]~FF .D_POLARITY = 1'b1;
    defparam \DESTINATION[2]~FF .SR_SYNC = 1'b1;
    defparam \DESTINATION[2]~FF .SR_VALUE = 1'b0;
    defparam \DESTINATION[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][0]~FF  (.D(n19664), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DESTINATION[1]~FF  (.D(\INSTRUCTION[16] ), .CE(n30664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DESTINATION[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \DESTINATION[1]~FF .CLK_POLARITY = 1'b1;
    defparam \DESTINATION[1]~FF .CE_POLARITY = 1'b1;
    defparam \DESTINATION[1]~FF .SR_POLARITY = 1'b1;
    defparam \DESTINATION[1]~FF .D_POLARITY = 1'b1;
    defparam \DESTINATION[1]~FF .SR_SYNC = 1'b1;
    defparam \DESTINATION[1]~FF .SR_VALUE = 1'b0;
    defparam \DESTINATION[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][0]~FF  (.D(n19664), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][0]~FF  (.D(n19664), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][0]~FF  (.D(n19664), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][0]~FF  (.D(n19664), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][0]~FF  (.D(n19664), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][0]~FF  (.D(n19664), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][0]~FF  (.D(n19664), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][0]~FF  (.D(n19664), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][0]~FF  (.D(n19664), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][0]~FF  (.D(n19664), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][0]~FF  (.D(n19664), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][0]~FF  (.D(n19664), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][0]~FF  (.D(n19664), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][0]~FF  (.D(n19664), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][0]~FF  (.D(n19664), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][0]~FF  (.D(n19664), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][0]~FF  (.D(n19664), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][0]~FF  (.D(n19664), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][0]~FF  (.D(n19664), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][0]~FF  (.D(n19664), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][0]~FF  (.D(n19664), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][0]~FF  (.D(n19664), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][0]~FF  (.D(n19664), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][0]~FF  (.D(n19664), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][0]~FF  (.D(n19664), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][0]~FF  (.D(n19664), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][0]~FF  (.D(n19664), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][0]~FF  (.D(n19664), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][0]~FF  (.D(n19664), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][0]~FF  (.D(n19664), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][0]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][0]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][0]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][0]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][0]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][0]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[20]~FF  (.D(n506_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[20]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[20]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[20]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[20]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[20]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[29]~FF  (.D(n497_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[29]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[29]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[29]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[29]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[29]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[28]~FF  (.D(n498_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[28]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[28]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[28]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[28]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[28]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ARG2[27]~FF  (.D(n499_2), .CE(n30664), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\ARG2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(544)
    defparam \ARG2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \ARG2[27]~FF .CE_POLARITY = 1'b1;
    defparam \ARG2[27]~FF .SR_POLARITY = 1'b1;
    defparam \ARG2[27]~FF .D_POLARITY = 1'b1;
    defparam \ARG2[27]~FF .SR_SYNC = 1'b1;
    defparam \ARG2[27]~FF .SR_VALUE = 1'b0;
    defparam \ARG2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[1]_2~FF  (.D(n1614), .CE(ceg_net408), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\RES[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \RES[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \RES[1]_2~FF .SR_POLARITY = 1'b1;
    defparam \RES[1]_2~FF .D_POLARITY = 1'b1;
    defparam \RES[1]_2~FF .SR_SYNC = 1'b1;
    defparam \RES[1]_2~FF .SR_VALUE = 1'b0;
    defparam \RES[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[2]_2~FF  (.D(n1613), .CE(ceg_net408), .CLK(\CLK~O ), .SR(1'b0), 
           .Q(\RES[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \RES[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \RES[2]_2~FF .SR_POLARITY = 1'b1;
    defparam \RES[2]_2~FF .D_POLARITY = 1'b1;
    defparam \RES[2]_2~FF .SR_SYNC = 1'b1;
    defparam \RES[2]_2~FF .SR_VALUE = 1'b0;
    defparam \RES[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i26  (.I0(n2756), .I1(1'b1), .CI(1'b0), 
            .CO(n5928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i27  (.I0(n2753), .I1(1'b1), .CI(1'b0), 
            .CO(n5927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i28  (.I0(n2750), .I1(1'b1), .CI(1'b0), 
            .CO(n5926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i29  (.I0(n2747), .I1(1'b1), .CI(1'b0), 
            .CO(n5925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i29 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i29 .I1_POLARITY = 1'b1;
    EFX_LUT4 \RES[15]_2~FF_brt_29_rtinv  (.I0(\RES[15]_2~FF_brt_29_q_pinv ), 
            .O(\RES[15]_2~FF_brt_29_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[15]_2~FF_brt_29_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[15]_2~FF_brt_30_brt_81  (.D(n5127), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[15]_2~FF_brt_30_brt_81_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[15]_2~FF_brt_30_brt_81 .CLK_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_81 .CE_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_81 .SR_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_81 .D_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_81 .SR_SYNC = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_81 .SR_VALUE = 1'b0;
    defparam \RES[15]_2~FF_brt_30_brt_81 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[9]_2~FF_brt_1_brt_24  (.D(n3547), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[9]_2~FF_brt_1_brt_24_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_1_brt_24 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_24 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_24 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_24 .D_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_24 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_24 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_24 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[9]_2~FF_brt_1_brt_23  (.D(n5039), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[9]_2~FF_brt_1_brt_23_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_1_brt_23 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_23 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_23 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_23 .D_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_23 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_23 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_23 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[7]_2~FF_brt_20_brt_70_brt_133_rtinv  (.I0(\RES[7]_2~FF_brt_20_brt_70_brt_133_q_pinv ), 
            .O(\RES[7]_2~FF_brt_20_brt_70_brt_133_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135  (.D(n1363), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135 .D_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_rtinv  (.I0(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_q_pinv ), 
            .O(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_rtinv .LUTMASK = 16'h5555;
    EFX_LUT4 \RES[22]_2~FF_brt_41_brt_98_rtinv  (.I0(\RES[22]_2~FF_brt_41_brt_98_q_pinv ), 
            .O(\RES[22]_2~FF_brt_41_brt_98_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[22]_2~FF_brt_41_brt_98_rtinv .LUTMASK = 16'h5555;
    EFX_LUT4 i17 (.I1(n221), .I2(RST), .I3(n1795), .O(n221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00FC */ ;
    defparam i17.LUTMASK = 16'h00FC;
    EFX_FF \RES[8]_2~FF_brt_22  (.D(n5037), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[8]_2~FF_brt_22_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[8]_2~FF_brt_22 .CLK_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_22 .CE_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_22 .SR_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_22 .D_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_22 .SR_SYNC = 1'b1;
    defparam \RES[8]_2~FF_brt_22 .SR_VALUE = 1'b0;
    defparam \RES[8]_2~FF_brt_22 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138  (.D(\OPERATION[0] ), 
           .CE(ceg_net408), .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138 .D_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[6]_2~FF_brt_131  (.D(n4999), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[6]_2~FF_brt_131_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[6]_2~FF_brt_131 .CLK_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_131 .CE_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_131 .SR_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_131 .D_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_131 .SR_SYNC = 1'b1;
    defparam \RES[6]_2~FF_brt_131 .SR_VALUE = 1'b0;
    defparam \RES[6]_2~FF_brt_131 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__4493 (.I0(STAGE2_EN), .I1(n51766), .O(n2953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4493.LUTMASK = 16'h8888;
    EFX_FF \RES[6]_2~FF_brt_130  (.D(n4997), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[6]_2~FF_brt_130_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[6]_2~FF_brt_130 .CLK_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_130 .CE_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_130 .SR_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_130 .D_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_130 .SR_SYNC = 1'b1;
    defparam \RES[6]_2~FF_brt_130 .SR_VALUE = 1'b0;
    defparam \RES[6]_2~FF_brt_130 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[6]_2~FF_brt_129  (.D(n4991), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[6]_2~FF_brt_129_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[6]_2~FF_brt_129 .CLK_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_129 .CE_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_129 .SR_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_129 .D_POLARITY = 1'b1;
    defparam \RES[6]_2~FF_brt_129 .SR_SYNC = 1'b1;
    defparam \RES[6]_2~FF_brt_129 .SR_VALUE = 1'b0;
    defparam \RES[6]_2~FF_brt_129 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[10]_2~FF_brt_3_brt_28_brt_75  (.D(n5058), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[10]_2~FF_brt_3_brt_28_brt_75_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_75 .CLK_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_75 .CE_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_75 .SR_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_75 .D_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_75 .SR_SYNC = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_75 .SR_VALUE = 1'b0;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_75 .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i32  (.I0(n2738), .I1(1'b1), .CI(1'b0), 
            .CO(n5922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i32 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i31  (.I0(n2741), .I1(1'b1), .CI(1'b0), 
            .CO(n5923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i31 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i31 .I1_POLARITY = 1'b1;
    EFX_FF \RES[4]_2~FF_brt_125  (.D(\OPERATION[3] ), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[4]_2~FF_brt_125_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[4]_2~FF_brt_125 .CLK_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_125 .CE_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_125 .SR_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_125 .D_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_125 .SR_SYNC = 1'b1;
    defparam \RES[4]_2~FF_brt_125 .SR_VALUE = 1'b0;
    defparam \RES[4]_2~FF_brt_125 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139  (.D(n1362), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139 .CLK_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139 .CE_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139 .SR_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139 .D_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139 .SR_SYNC = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139 .SR_VALUE = 1'b0;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[8]_2~FF_brt_21_brt_71  (.D(n5026), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[8]_2~FF_brt_21_brt_71_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[8]_2~FF_brt_21_brt_71 .CLK_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_71 .CE_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_71 .SR_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_71 .D_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_71 .SR_SYNC = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_71 .SR_VALUE = 1'b0;
    defparam \RES[8]_2~FF_brt_21_brt_71 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[7]_2~FF_brt_19  (.D(n5000), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[7]_2~FF_brt_19_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[7]_2~FF_brt_19 .CLK_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_19 .CE_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_19 .SR_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_19 .D_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_19 .SR_SYNC = 1'b1;
    defparam \RES[7]_2~FF_brt_19 .SR_VALUE = 1'b0;
    defparam \RES[7]_2~FF_brt_19 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[7]_2~FF_brt_18  (.D(n5004), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[7]_2~FF_brt_18_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[7]_2~FF_brt_18 .CLK_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_18 .CE_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_18 .SR_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_18 .D_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_18 .SR_SYNC = 1'b1;
    defparam \RES[7]_2~FF_brt_18 .SR_VALUE = 1'b0;
    defparam \RES[7]_2~FF_brt_18 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[0]_2~FF_brt_193  (.D(n3551), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[0]_2~FF_brt_193_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[0]_2~FF_brt_193 .CLK_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_193 .CE_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_193 .SR_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_193 .D_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_193 .SR_SYNC = 1'b1;
    defparam \RES[0]_2~FF_brt_193 .SR_VALUE = 1'b0;
    defparam \RES[0]_2~FF_brt_193 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[7]_2~FF_brt_20_brt_68  (.D(n5016), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[7]_2~FF_brt_20_brt_68_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[7]_2~FF_brt_20_brt_68 .CLK_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_68 .CE_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_68 .SR_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_68 .D_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_68 .SR_SYNC = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_68 .SR_VALUE = 1'b0;
    defparam \RES[7]_2~FF_brt_20_brt_68 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \GPR[1]~FF  (.D(\DESTINATION[1] ), .CE(n30678), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\GPR[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \GPR[1]~FF .CLK_POLARITY = 1'b1;
    defparam \GPR[1]~FF .CE_POLARITY = 1'b1;
    defparam \GPR[1]~FF .SR_POLARITY = 1'b1;
    defparam \GPR[1]~FF .D_POLARITY = 1'b1;
    defparam \GPR[1]~FF .SR_SYNC = 1'b1;
    defparam \GPR[1]~FF .SR_VALUE = 1'b0;
    defparam \GPR[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \GPR[2]~FF  (.D(\DESTINATION[2] ), .CE(n30678), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\GPR[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \GPR[2]~FF .CLK_POLARITY = 1'b1;
    defparam \GPR[2]~FF .CE_POLARITY = 1'b1;
    defparam \GPR[2]~FF .SR_POLARITY = 1'b1;
    defparam \GPR[2]~FF .D_POLARITY = 1'b1;
    defparam \GPR[2]~FF .SR_SYNC = 1'b1;
    defparam \GPR[2]~FF .SR_VALUE = 1'b0;
    defparam \GPR[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \GPR[3]~FF  (.D(\DESTINATION[3] ), .CE(n30678), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\GPR[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \GPR[3]~FF .CLK_POLARITY = 1'b1;
    defparam \GPR[3]~FF .CE_POLARITY = 1'b1;
    defparam \GPR[3]~FF .SR_POLARITY = 1'b1;
    defparam \GPR[3]~FF .D_POLARITY = 1'b1;
    defparam \GPR[3]~FF .SR_SYNC = 1'b1;
    defparam \GPR[3]~FF .SR_VALUE = 1'b0;
    defparam \GPR[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \GPR[4]~FF  (.D(\DESTINATION[4] ), .CE(n30678), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\GPR[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \GPR[4]~FF .CLK_POLARITY = 1'b1;
    defparam \GPR[4]~FF .CE_POLARITY = 1'b1;
    defparam \GPR[4]~FF .SR_POLARITY = 1'b1;
    defparam \GPR[4]~FF .D_POLARITY = 1'b1;
    defparam \GPR[4]~FF .SR_SYNC = 1'b1;
    defparam \GPR[4]~FF .SR_VALUE = 1'b0;
    defparam \GPR[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DATA_FORMAT_2[1]~FF  (.D(\DATA_FORMAT[1] ), .CE(n50476), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DATA_FORMAT_2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \DATA_FORMAT_2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[1]~FF .CE_POLARITY = 1'b0;
    defparam \DATA_FORMAT_2[1]~FF .SR_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[1]~FF .D_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[1]~FF .SR_SYNC = 1'b1;
    defparam \DATA_FORMAT_2[1]~FF .SR_VALUE = 1'b0;
    defparam \DATA_FORMAT_2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DATA_FORMAT_2[2]~FF  (.D(\DATA_FORMAT[2] ), .CE(n50476), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\DATA_FORMAT_2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \DATA_FORMAT_2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[2]~FF .CE_POLARITY = 1'b0;
    defparam \DATA_FORMAT_2[2]~FF .SR_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[2]~FF .D_POLARITY = 1'b1;
    defparam \DATA_FORMAT_2[2]~FF .SR_SYNC = 1'b1;
    defparam \DATA_FORMAT_2[2]~FF .SR_VALUE = 1'b0;
    defparam \DATA_FORMAT_2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[1]~FF  (.D(n1387), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[1]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[1]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[1]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[1]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[1]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[1]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[2]~FF  (.D(n1385), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[2]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[2]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[2]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[2]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[2]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[2]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[3]~FF  (.D(n1383), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[3]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[3]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[3]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[3]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[3]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[3]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[4]~FF  (.D(n1381), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[4]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[4]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[4]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[4]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[4]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[4]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[5]~FF  (.D(n1379), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[5]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[5]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[5]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[5]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[5]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[5]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[6]~FF  (.D(n1377), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[6]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[6]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[6]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[6]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[6]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[6]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[7]~FF  (.D(n1375), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[7]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[7]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[7]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[7]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[7]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[7]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[8]~FF  (.D(n1373), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[8]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[8]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[8]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[8]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[8]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[8]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_ADDRESS[9]~FF  (.D(n1372), .CE(n50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_ADDRESS[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_ADDRESS[9]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[9]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[9]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[9]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_ADDRESS[9]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_ADDRESS[9]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_ADDRESS[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[1]~FF  (.D(\ARG2[1] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[1]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[1]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[1]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[1]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[1]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[2]~FF  (.D(\ARG2[2] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[2]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[2]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[2]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[2]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[2]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[3]~FF  (.D(\ARG2[3] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[3]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[3]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[3]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[3]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[3]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[4]~FF  (.D(\ARG2[4] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[4]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[4]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[4]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[4]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[4]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[5]~FF  (.D(\ARG2[5] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[5]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[5]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[5]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[5]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[5]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[6]~FF  (.D(\ARG2[6] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[6]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[6]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[6]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[6]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[6]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[7]~FF  (.D(\ARG2[7] ), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[7]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[7]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[7]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[7]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[7]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[8]~FF  (.D(n1575), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[8]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[8]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[8]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[8]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[8]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[9]~FF  (.D(n1574_2), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[9]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[9]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[9]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[9]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[9]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[9]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[10]~FF  (.D(n1573), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[10]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[10]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[10]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[10]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[10]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[10]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[11]~FF  (.D(n1572), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[11]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[11]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[11]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[11]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[11]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[11]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[12]~FF  (.D(n1571), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[12]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[12]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[12]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[12]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[12]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[12]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[13]~FF  (.D(n1570), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[13]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[13]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[13]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[13]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[13]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[13]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[14]~FF  (.D(n1569), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[14]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[14]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[14]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[14]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[14]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[14]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[15]~FF  (.D(n1568), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[15]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[15]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[15]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[15]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[15]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[15]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[16]~FF  (.D(n1567), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[16]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[16]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[16]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[16]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[16]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[16]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[17]~FF  (.D(n1566), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[17]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[17]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[17]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[17]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[17]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[17]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[18]~FF  (.D(n1565), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[18]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[18]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[18]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[18]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[18]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[18]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[19]~FF  (.D(n1564), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[19]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[19]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[19]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[19]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[19]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[19]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[20]~FF  (.D(n1563), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[20]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[20]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[20]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[20]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[20]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[20]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[21]~FF  (.D(n1562), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[21]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[21]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[21]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[21]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[21]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[21]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[22]~FF  (.D(n1561), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[22]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[22]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[22]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[22]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[22]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[22]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[23]~FF  (.D(n1560), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[23]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[23]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[23]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[23]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[23]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[23]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[24]~FF  (.D(n1559), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[24]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[24]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[24]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[24]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[24]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[24]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[25]~FF  (.D(n1558), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[25]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[25]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[25]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[25]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[25]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[25]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[26]~FF  (.D(n1557), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[26]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[26]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[26]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[26]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[26]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[26]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[27]~FF  (.D(n1556), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[27]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[27]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[27]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[27]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[27]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[27]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[28]~FF  (.D(n1555), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[28]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[28]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[28]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[28]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[28]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[28]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[29]~FF  (.D(n1554), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[29]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[29]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[29]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[29]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[29]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[29]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[30]~FF  (.D(n1553), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[30]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[30]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[30]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[30]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[30]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[30]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \SAVE_DATA[31]~FF  (.D(n1552), .CE(ceg_net35302), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\SAVE_DATA[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \SAVE_DATA[31]~FF .CLK_POLARITY = 1'b1;
    defparam \SAVE_DATA[31]~FF .CE_POLARITY = 1'b1;
    defparam \SAVE_DATA[31]~FF .SR_POLARITY = 1'b1;
    defparam \SAVE_DATA[31]~FF .D_POLARITY = 1'b1;
    defparam \SAVE_DATA[31]~FF .SR_SYNC = 1'b1;
    defparam \SAVE_DATA[31]~FF .SR_VALUE = 1'b0;
    defparam \SAVE_DATA[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][8]~FF  (.D(n17577), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][9]~FF  (.D(n17576), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][10]~FF  (.D(n17575), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][11]~FF  (.D(n17574), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][12]~FF  (.D(n17573), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][13]~FF  (.D(n17572), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][14]~FF  (.D(n17571), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][15]~FF  (.D(n17570), .CE(ceg_net41512), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][16]~FF  (.D(n17569), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][17]~FF  (.D(n17568), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][18]~FF  (.D(n17567), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][19]~FF  (.D(n17566), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][20]~FF  (.D(n17565), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][21]~FF  (.D(n17564), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][22]~FF  (.D(n17563), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][23]~FF  (.D(n17562), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][24]~FF  (.D(n17561), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][25]~FF  (.D(n17560), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][26]~FF  (.D(n17559), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][27]~FF  (.D(n17558), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][28]~FF  (.D(n17557), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][29]~FF  (.D(n17556), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][30]~FF  (.D(n17555), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[0][31]~FF  (.D(n17554), .CE(ceg_net49709), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[0][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[0][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[0][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[0][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[0][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[0][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[0][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[0][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][8]~FF  (.D(n17610), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][9]~FF  (.D(n17609), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][10]~FF  (.D(n17608), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][11]~FF  (.D(n17607), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][12]~FF  (.D(n17606), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][13]~FF  (.D(n17605), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][14]~FF  (.D(n17604), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][15]~FF  (.D(n17603), .CE(ceg_net41704), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][16]~FF  (.D(n17602), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][17]~FF  (.D(n17601), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][18]~FF  (.D(n17600), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][19]~FF  (.D(n17599), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][20]~FF  (.D(n17598), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][21]~FF  (.D(n17597), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][22]~FF  (.D(n17596), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][23]~FF  (.D(n17595), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][24]~FF  (.D(n17594), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][25]~FF  (.D(n17593), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][26]~FF  (.D(n17592), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][27]~FF  (.D(n17591), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][28]~FF  (.D(n17590), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][29]~FF  (.D(n17589), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][30]~FF  (.D(n17588), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[1][31]~FF  (.D(n17587), .CE(ceg_net49773), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[1][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[1][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[1][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[1][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[1][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[1][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[1][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[1][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][8]~FF  (.D(n17643), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][9]~FF  (.D(n17642), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][10]~FF  (.D(n17641), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][11]~FF  (.D(n17640), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][12]~FF  (.D(n17639), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][13]~FF  (.D(n17638), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][14]~FF  (.D(n17637), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][15]~FF  (.D(n17636), .CE(ceg_net41896), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][16]~FF  (.D(n17635), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][17]~FF  (.D(n17634), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][18]~FF  (.D(n17633), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][19]~FF  (.D(n17632), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][20]~FF  (.D(n17631), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][21]~FF  (.D(n17630), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][22]~FF  (.D(n17629), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][23]~FF  (.D(n17628), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][24]~FF  (.D(n17627), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][25]~FF  (.D(n17626), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][26]~FF  (.D(n17625), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][27]~FF  (.D(n17624), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][28]~FF  (.D(n17623), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][29]~FF  (.D(n17622), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][30]~FF  (.D(n17621), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[2][31]~FF  (.D(n17620), .CE(ceg_net49837), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[2][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[2][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[2][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[2][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[2][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[2][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[2][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[2][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][8]~FF  (.D(n17676), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][9]~FF  (.D(n17675), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][10]~FF  (.D(n17674), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][11]~FF  (.D(n17673), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][12]~FF  (.D(n17672), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][13]~FF  (.D(n17671), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][14]~FF  (.D(n17670), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][15]~FF  (.D(n17669), .CE(ceg_net42088), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][16]~FF  (.D(n17668), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][17]~FF  (.D(n17667), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][18]~FF  (.D(n17666), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][19]~FF  (.D(n17665), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][20]~FF  (.D(n17664), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][21]~FF  (.D(n17663), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][22]~FF  (.D(n17662), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][23]~FF  (.D(n17661), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][24]~FF  (.D(n17660), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][25]~FF  (.D(n17659), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][26]~FF  (.D(n17658), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][27]~FF  (.D(n17657), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][28]~FF  (.D(n17656), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][29]~FF  (.D(n17655), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][30]~FF  (.D(n17654), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[3][31]~FF  (.D(n17653), .CE(ceg_net49901), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[3][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[3][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[3][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[3][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[3][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[3][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[3][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[3][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][8]~FF  (.D(n17709), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][9]~FF  (.D(n17708), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][10]~FF  (.D(n17707), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][11]~FF  (.D(n17706), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][12]~FF  (.D(n17705), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][13]~FF  (.D(n17704), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][14]~FF  (.D(n17703), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][15]~FF  (.D(n17702), .CE(ceg_net42280), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][16]~FF  (.D(n17701), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][17]~FF  (.D(n17700), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][18]~FF  (.D(n17699), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][19]~FF  (.D(n17698), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][20]~FF  (.D(n17697), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][21]~FF  (.D(n17696), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][22]~FF  (.D(n17695), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][23]~FF  (.D(n17694), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][24]~FF  (.D(n17693), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][25]~FF  (.D(n17692), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][26]~FF  (.D(n17691), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][27]~FF  (.D(n17690), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][28]~FF  (.D(n17689), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][29]~FF  (.D(n17688), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][30]~FF  (.D(n17687), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[4][31]~FF  (.D(n17686), .CE(ceg_net49965), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[4][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[4][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[4][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[4][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[4][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[4][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[4][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[4][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][8]~FF  (.D(n17742), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][9]~FF  (.D(n17741), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][10]~FF  (.D(n17740), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][11]~FF  (.D(n17739), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][12]~FF  (.D(n17738), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][13]~FF  (.D(n17737), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][14]~FF  (.D(n17736), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][15]~FF  (.D(n17735), .CE(ceg_net42472), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][16]~FF  (.D(n17734), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][17]~FF  (.D(n17733), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][18]~FF  (.D(n17732), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][19]~FF  (.D(n17731), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][20]~FF  (.D(n17730), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][21]~FF  (.D(n17729), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][22]~FF  (.D(n17728), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][23]~FF  (.D(n17727), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][24]~FF  (.D(n17726), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][25]~FF  (.D(n17725), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][26]~FF  (.D(n17724), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][27]~FF  (.D(n17723), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][28]~FF  (.D(n17722), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][29]~FF  (.D(n17721), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][30]~FF  (.D(n17720), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[5][31]~FF  (.D(n17719), .CE(ceg_net50029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[5][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[5][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[5][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[5][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[5][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[5][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[5][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[5][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][8]~FF  (.D(n17775), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][9]~FF  (.D(n17774), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][10]~FF  (.D(n17773), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][11]~FF  (.D(n17772), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][12]~FF  (.D(n17771), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][13]~FF  (.D(n17770), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][14]~FF  (.D(n17769), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][15]~FF  (.D(n17768), .CE(ceg_net42664), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][16]~FF  (.D(n17767), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][17]~FF  (.D(n17766), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][18]~FF  (.D(n17765), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][19]~FF  (.D(n17764), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][20]~FF  (.D(n17763), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][21]~FF  (.D(n17762), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][22]~FF  (.D(n17761), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][23]~FF  (.D(n17760), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][24]~FF  (.D(n17759), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][25]~FF  (.D(n17758), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][26]~FF  (.D(n17757), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][27]~FF  (.D(n17756), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][28]~FF  (.D(n17755), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][29]~FF  (.D(n17754), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][30]~FF  (.D(n17753), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[6][31]~FF  (.D(n17752), .CE(ceg_net50093), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[6][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[6][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[6][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[6][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[6][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[6][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[6][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[6][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][8]~FF  (.D(n17808), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][9]~FF  (.D(n17807), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][10]~FF  (.D(n17806), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][11]~FF  (.D(n17805), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][12]~FF  (.D(n17804), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][13]~FF  (.D(n17803), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][14]~FF  (.D(n17802), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][15]~FF  (.D(n17801), .CE(ceg_net42856), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][16]~FF  (.D(n17800), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][17]~FF  (.D(n17799), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][18]~FF  (.D(n17798), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][19]~FF  (.D(n17797), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][20]~FF  (.D(n17796), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][21]~FF  (.D(n17795), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][22]~FF  (.D(n17794), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][23]~FF  (.D(n17793), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][24]~FF  (.D(n17792), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][25]~FF  (.D(n17791), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][26]~FF  (.D(n17790), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][27]~FF  (.D(n17789), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][28]~FF  (.D(n17788), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][29]~FF  (.D(n17787), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][30]~FF  (.D(n17786), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[7][31]~FF  (.D(n17785), .CE(ceg_net50157), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[7][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[7][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[7][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[7][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[7][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[7][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[7][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[7][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][8]~FF  (.D(n17841), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][9]~FF  (.D(n17840), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][10]~FF  (.D(n17839), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][11]~FF  (.D(n17838), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][12]~FF  (.D(n17837), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][13]~FF  (.D(n17836), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][14]~FF  (.D(n17835), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][15]~FF  (.D(n17834), .CE(ceg_net43048), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][16]~FF  (.D(n17833), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][17]~FF  (.D(n17832), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][18]~FF  (.D(n17831), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][19]~FF  (.D(n17830), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][20]~FF  (.D(n17829), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][21]~FF  (.D(n17828), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][22]~FF  (.D(n17827), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][23]~FF  (.D(n17826), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][24]~FF  (.D(n17825), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][25]~FF  (.D(n17824), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][26]~FF  (.D(n17823), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][27]~FF  (.D(n17822), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][28]~FF  (.D(n17821), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][29]~FF  (.D(n17820), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][30]~FF  (.D(n17819), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[8][31]~FF  (.D(n17818), .CE(ceg_net50221), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[8][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[8][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[8][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[8][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[8][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[8][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[8][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[8][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][8]~FF  (.D(n17874), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][9]~FF  (.D(n17873), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][10]~FF  (.D(n17872), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][11]~FF  (.D(n17871), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][12]~FF  (.D(n17870), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][13]~FF  (.D(n17869), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][14]~FF  (.D(n17868), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][15]~FF  (.D(n17867), .CE(ceg_net43240), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][16]~FF  (.D(n17866), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][17]~FF  (.D(n17865), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][18]~FF  (.D(n17864), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][19]~FF  (.D(n17863), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][20]~FF  (.D(n17862), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][21]~FF  (.D(n17861), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][22]~FF  (.D(n17860), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][23]~FF  (.D(n17859), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][24]~FF  (.D(n17858), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][25]~FF  (.D(n17857), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][26]~FF  (.D(n17856), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][27]~FF  (.D(n17855), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][28]~FF  (.D(n17854), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][29]~FF  (.D(n17853), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][30]~FF  (.D(n17852), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[9][31]~FF  (.D(n17851), .CE(ceg_net50285), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[9][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[9][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[9][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[9][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[9][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[9][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[9][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[9][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][8]~FF  (.D(n17907), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][9]~FF  (.D(n17906), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][10]~FF  (.D(n17905), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][11]~FF  (.D(n17904), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][12]~FF  (.D(n17903), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][13]~FF  (.D(n17902), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][14]~FF  (.D(n17901), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][15]~FF  (.D(n17900), .CE(ceg_net43432), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][16]~FF  (.D(n17899), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][17]~FF  (.D(n17898), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][18]~FF  (.D(n17897), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][19]~FF  (.D(n17896), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][20]~FF  (.D(n17895), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][21]~FF  (.D(n17894), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][22]~FF  (.D(n17893), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][23]~FF  (.D(n17892), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][24]~FF  (.D(n17891), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][25]~FF  (.D(n17890), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][26]~FF  (.D(n17889), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][27]~FF  (.D(n17888), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][28]~FF  (.D(n17887), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][29]~FF  (.D(n17886), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][30]~FF  (.D(n17885), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[10][31]~FF  (.D(n17884), .CE(ceg_net50349), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[10][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[10][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[10][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[10][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[10][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[10][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[10][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[10][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][8]~FF  (.D(n17940), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][9]~FF  (.D(n17939), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][10]~FF  (.D(n17938), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][11]~FF  (.D(n17937), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][12]~FF  (.D(n17936), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][13]~FF  (.D(n17935), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][14]~FF  (.D(n17934), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][15]~FF  (.D(n17933), .CE(ceg_net43624), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][16]~FF  (.D(n17932), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][17]~FF  (.D(n17931), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][18]~FF  (.D(n17930), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][19]~FF  (.D(n17929), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][20]~FF  (.D(n17928), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][21]~FF  (.D(n17927), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][22]~FF  (.D(n17926), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][23]~FF  (.D(n17925), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][24]~FF  (.D(n17924), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][25]~FF  (.D(n17923), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][26]~FF  (.D(n17922), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][27]~FF  (.D(n17921), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][28]~FF  (.D(n17920), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][29]~FF  (.D(n17919), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][30]~FF  (.D(n17918), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[11][31]~FF  (.D(n17917), .CE(ceg_net50413), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[11][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[11][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[11][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[11][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[11][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[11][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[11][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[11][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][8]~FF  (.D(n17973), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][9]~FF  (.D(n17972), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][10]~FF  (.D(n17971), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][11]~FF  (.D(n17970), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][12]~FF  (.D(n17969), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][13]~FF  (.D(n17968), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][14]~FF  (.D(n17967), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][15]~FF  (.D(n17966), .CE(ceg_net43816), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][16]~FF  (.D(n17965), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][17]~FF  (.D(n17964), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][18]~FF  (.D(n17963), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][19]~FF  (.D(n17962), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][20]~FF  (.D(n17961), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][21]~FF  (.D(n17960), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][22]~FF  (.D(n17959), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][23]~FF  (.D(n17958), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][24]~FF  (.D(n17957), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][25]~FF  (.D(n17956), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][26]~FF  (.D(n17955), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][27]~FF  (.D(n17954), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][28]~FF  (.D(n17953), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][29]~FF  (.D(n17952), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][30]~FF  (.D(n17951), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[12][31]~FF  (.D(n17950), .CE(ceg_net50477), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[12][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[12][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[12][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[12][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[12][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[12][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[12][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[12][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][8]~FF  (.D(n18006), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][9]~FF  (.D(n18005), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][10]~FF  (.D(n18004), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][11]~FF  (.D(n18003), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][12]~FF  (.D(n18002), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][13]~FF  (.D(n18001), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][14]~FF  (.D(n18000), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][15]~FF  (.D(n17999), .CE(ceg_net44008), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][16]~FF  (.D(n17998), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][17]~FF  (.D(n17997), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][18]~FF  (.D(n17996), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][19]~FF  (.D(n17995), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][20]~FF  (.D(n17994), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][21]~FF  (.D(n17993), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][22]~FF  (.D(n17992), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][23]~FF  (.D(n17991), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][24]~FF  (.D(n17990), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][25]~FF  (.D(n17989), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][26]~FF  (.D(n17988), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][27]~FF  (.D(n17987), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][28]~FF  (.D(n17986), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][29]~FF  (.D(n17985), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][30]~FF  (.D(n17984), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[13][31]~FF  (.D(n17983), .CE(ceg_net50541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[13][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[13][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[13][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[13][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[13][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[13][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[13][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[13][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][8]~FF  (.D(n18039), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][9]~FF  (.D(n18038), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][10]~FF  (.D(n18037), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][11]~FF  (.D(n18036), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][12]~FF  (.D(n18035), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][13]~FF  (.D(n18034), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][14]~FF  (.D(n18033), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][15]~FF  (.D(n18032), .CE(ceg_net44200), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][16]~FF  (.D(n18031), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][17]~FF  (.D(n18030), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][18]~FF  (.D(n18029), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][19]~FF  (.D(n18028), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][20]~FF  (.D(n18027), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][21]~FF  (.D(n18026), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][22]~FF  (.D(n18025), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][23]~FF  (.D(n18024), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][24]~FF  (.D(n18023), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][25]~FF  (.D(n18022), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][26]~FF  (.D(n18021), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][27]~FF  (.D(n18020), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][28]~FF  (.D(n18019), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][29]~FF  (.D(n18018), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][30]~FF  (.D(n18017), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[14][31]~FF  (.D(n18016), .CE(ceg_net50605), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[14][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[14][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[14][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[14][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[14][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[14][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[14][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[14][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][8]~FF  (.D(n18072), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][9]~FF  (.D(n18071), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][10]~FF  (.D(n18070), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][11]~FF  (.D(n18069), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][12]~FF  (.D(n18068), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][13]~FF  (.D(n18067), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][14]~FF  (.D(n18066), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][15]~FF  (.D(n18065), .CE(ceg_net44392), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][16]~FF  (.D(n18064), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][17]~FF  (.D(n18063), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][18]~FF  (.D(n18062), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][19]~FF  (.D(n18061), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][20]~FF  (.D(n18060), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][21]~FF  (.D(n18059), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][22]~FF  (.D(n18058), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][23]~FF  (.D(n18057), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][24]~FF  (.D(n18056), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][25]~FF  (.D(n18055), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][26]~FF  (.D(n18054), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][27]~FF  (.D(n18053), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][28]~FF  (.D(n18052), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][29]~FF  (.D(n18051), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][30]~FF  (.D(n18050), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[15][31]~FF  (.D(n18049), .CE(ceg_net50669), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[15][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[15][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[15][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[15][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[15][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[15][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[15][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[15][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][8]~FF  (.D(n18105), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][9]~FF  (.D(n18104), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][10]~FF  (.D(n18103), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][11]~FF  (.D(n18102), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][12]~FF  (.D(n18101), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][13]~FF  (.D(n18100), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][14]~FF  (.D(n18099), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][15]~FF  (.D(n18098), .CE(ceg_net44584), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][16]~FF  (.D(n18097), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][17]~FF  (.D(n18096), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][18]~FF  (.D(n18095), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][19]~FF  (.D(n18094), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][20]~FF  (.D(n18093), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][21]~FF  (.D(n18092), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][22]~FF  (.D(n18091), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][23]~FF  (.D(n18090), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][24]~FF  (.D(n18089), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][25]~FF  (.D(n18088), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][26]~FF  (.D(n18087), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][27]~FF  (.D(n18086), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][28]~FF  (.D(n18085), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][29]~FF  (.D(n18084), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][30]~FF  (.D(n18083), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[16][31]~FF  (.D(n18082), .CE(ceg_net50733), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[16][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[16][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[16][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[16][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[16][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[16][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[16][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[16][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][8]~FF  (.D(n18138), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][9]~FF  (.D(n18137), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][10]~FF  (.D(n18136), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][11]~FF  (.D(n18135), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][12]~FF  (.D(n18134), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][13]~FF  (.D(n18133), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][14]~FF  (.D(n18132), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][15]~FF  (.D(n18131), .CE(ceg_net44776), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][16]~FF  (.D(n18130), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][17]~FF  (.D(n18129), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][18]~FF  (.D(n18128), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][19]~FF  (.D(n18127), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][20]~FF  (.D(n18126), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][21]~FF  (.D(n18125), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][22]~FF  (.D(n18124), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][23]~FF  (.D(n18123), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][24]~FF  (.D(n18122), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][25]~FF  (.D(n18121), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][26]~FF  (.D(n18120), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][27]~FF  (.D(n18119), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][28]~FF  (.D(n18118), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][29]~FF  (.D(n18117), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][30]~FF  (.D(n18116), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[17][31]~FF  (.D(n18115), .CE(ceg_net50797), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[17][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[17][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[17][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[17][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[17][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[17][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[17][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[17][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][8]~FF  (.D(n18171), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][9]~FF  (.D(n18170), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][10]~FF  (.D(n18169), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][11]~FF  (.D(n18168), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][12]~FF  (.D(n18167), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][13]~FF  (.D(n18166), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][14]~FF  (.D(n18165), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][15]~FF  (.D(n18164), .CE(ceg_net44968), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][16]~FF  (.D(n18163), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][17]~FF  (.D(n18162), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][18]~FF  (.D(n18161), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][19]~FF  (.D(n18160), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][20]~FF  (.D(n18159), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][21]~FF  (.D(n18158), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][22]~FF  (.D(n18157), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][23]~FF  (.D(n18156), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][24]~FF  (.D(n18155), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][25]~FF  (.D(n18154), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][26]~FF  (.D(n18153), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][27]~FF  (.D(n18152), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][28]~FF  (.D(n18151), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][29]~FF  (.D(n18150), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][30]~FF  (.D(n18149), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[18][31]~FF  (.D(n18148), .CE(ceg_net50861), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[18][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[18][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[18][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[18][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[18][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[18][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[18][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[18][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][8]~FF  (.D(n18204), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][9]~FF  (.D(n18203), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][10]~FF  (.D(n18202), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][11]~FF  (.D(n18201), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][12]~FF  (.D(n18200), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][13]~FF  (.D(n18199), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][14]~FF  (.D(n18198), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][15]~FF  (.D(n18197), .CE(ceg_net45160), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][16]~FF  (.D(n18196), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][17]~FF  (.D(n18195), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][18]~FF  (.D(n18194), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][19]~FF  (.D(n18193), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][20]~FF  (.D(n18192), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][21]~FF  (.D(n18191), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][22]~FF  (.D(n18190), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][23]~FF  (.D(n18189), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][24]~FF  (.D(n18188), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][25]~FF  (.D(n18187), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][26]~FF  (.D(n18186), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][27]~FF  (.D(n18185), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][28]~FF  (.D(n18184), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][29]~FF  (.D(n18183), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][30]~FF  (.D(n18182), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[19][31]~FF  (.D(n18181), .CE(ceg_net50925), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[19][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[19][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[19][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[19][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[19][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[19][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[19][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[19][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][8]~FF  (.D(n18237), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][9]~FF  (.D(n18236), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][10]~FF  (.D(n18235), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][11]~FF  (.D(n18234), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][12]~FF  (.D(n18233), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][13]~FF  (.D(n18232), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][14]~FF  (.D(n18231), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][15]~FF  (.D(n18230), .CE(ceg_net45352), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][16]~FF  (.D(n18229), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][17]~FF  (.D(n18228), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][18]~FF  (.D(n18227), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][19]~FF  (.D(n18226), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][20]~FF  (.D(n18225), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][21]~FF  (.D(n18224), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][22]~FF  (.D(n18223), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][23]~FF  (.D(n18222), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][24]~FF  (.D(n18221), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][25]~FF  (.D(n18220), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][26]~FF  (.D(n18219), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][27]~FF  (.D(n18218), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][28]~FF  (.D(n18217), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][29]~FF  (.D(n18216), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][30]~FF  (.D(n18215), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[20][31]~FF  (.D(n18214), .CE(ceg_net50989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[20][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[20][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[20][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[20][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[20][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[20][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[20][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[20][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][8]~FF  (.D(n18270), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][9]~FF  (.D(n18269), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][10]~FF  (.D(n18268), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][11]~FF  (.D(n18267), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][12]~FF  (.D(n18266), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][13]~FF  (.D(n18265), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][14]~FF  (.D(n18264), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][15]~FF  (.D(n18263), .CE(ceg_net45544), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][16]~FF  (.D(n18262), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][17]~FF  (.D(n18261), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][18]~FF  (.D(n18260), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][19]~FF  (.D(n18259), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][20]~FF  (.D(n18258), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][21]~FF  (.D(n18257), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][22]~FF  (.D(n18256), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][23]~FF  (.D(n18255), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][24]~FF  (.D(n18254), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][25]~FF  (.D(n18253), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][26]~FF  (.D(n18252), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][27]~FF  (.D(n18251), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][28]~FF  (.D(n18250), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][29]~FF  (.D(n18249), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][30]~FF  (.D(n18248), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[21][31]~FF  (.D(n18247), .CE(ceg_net51053), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[21][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[21][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[21][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[21][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[21][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[21][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[21][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[21][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][8]~FF  (.D(n18303), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][9]~FF  (.D(n18302), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][10]~FF  (.D(n18301), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][11]~FF  (.D(n18300), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][12]~FF  (.D(n18299), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][13]~FF  (.D(n18298), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][14]~FF  (.D(n18297), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][15]~FF  (.D(n18296), .CE(ceg_net45736), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][16]~FF  (.D(n18295), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][17]~FF  (.D(n18294), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][18]~FF  (.D(n18293), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][19]~FF  (.D(n18292), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][20]~FF  (.D(n18291), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][21]~FF  (.D(n18290), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][22]~FF  (.D(n18289), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][23]~FF  (.D(n18288), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][24]~FF  (.D(n18287), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][25]~FF  (.D(n18286), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][26]~FF  (.D(n18285), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][27]~FF  (.D(n18284), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][28]~FF  (.D(n18283), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][29]~FF  (.D(n18282), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][30]~FF  (.D(n18281), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[22][31]~FF  (.D(n18280), .CE(ceg_net51117), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[22][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[22][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[22][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[22][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[22][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[22][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[22][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[22][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][8]~FF  (.D(n18336), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][9]~FF  (.D(n18335), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][10]~FF  (.D(n18334), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][11]~FF  (.D(n18333), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][12]~FF  (.D(n18332), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][13]~FF  (.D(n18331), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][14]~FF  (.D(n18330), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][15]~FF  (.D(n18329), .CE(ceg_net45928), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][16]~FF  (.D(n18328), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][17]~FF  (.D(n18327), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][18]~FF  (.D(n18326), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][19]~FF  (.D(n18325), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][20]~FF  (.D(n18324), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][21]~FF  (.D(n18323), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][22]~FF  (.D(n18322), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][23]~FF  (.D(n18321), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][24]~FF  (.D(n18320), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][25]~FF  (.D(n18319), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][26]~FF  (.D(n18318), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][27]~FF  (.D(n18317), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][28]~FF  (.D(n18316), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][29]~FF  (.D(n18315), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][30]~FF  (.D(n18314), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[23][31]~FF  (.D(n18313), .CE(ceg_net51181), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[23][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[23][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[23][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[23][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[23][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[23][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[23][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[23][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][8]~FF  (.D(n18369), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][9]~FF  (.D(n18368), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][10]~FF  (.D(n18367), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][11]~FF  (.D(n18366), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][12]~FF  (.D(n18365), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][13]~FF  (.D(n18364), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][14]~FF  (.D(n18363), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][15]~FF  (.D(n18362), .CE(ceg_net46120), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][16]~FF  (.D(n18361), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][17]~FF  (.D(n18360), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][18]~FF  (.D(n18359), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][19]~FF  (.D(n18358), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][20]~FF  (.D(n18357), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][21]~FF  (.D(n18356), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][22]~FF  (.D(n18355), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][23]~FF  (.D(n18354), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][24]~FF  (.D(n18353), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][25]~FF  (.D(n18352), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][26]~FF  (.D(n18351), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][27]~FF  (.D(n18350), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][28]~FF  (.D(n18349), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][29]~FF  (.D(n18348), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][30]~FF  (.D(n18347), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[24][31]~FF  (.D(n18346), .CE(ceg_net51245), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[24][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[24][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[24][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[24][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[24][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[24][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[24][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[24][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][8]~FF  (.D(n18402), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][9]~FF  (.D(n18401), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][10]~FF  (.D(n18400), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][11]~FF  (.D(n18399), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][12]~FF  (.D(n18398), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][13]~FF  (.D(n18397), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][14]~FF  (.D(n18396), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][15]~FF  (.D(n18395), .CE(ceg_net46312), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][16]~FF  (.D(n18394), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][17]~FF  (.D(n18393), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][18]~FF  (.D(n18392), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][19]~FF  (.D(n18391), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][20]~FF  (.D(n18390), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][21]~FF  (.D(n18389), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][22]~FF  (.D(n18388), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][23]~FF  (.D(n18387), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][24]~FF  (.D(n18386), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][25]~FF  (.D(n18385), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][26]~FF  (.D(n18384), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][27]~FF  (.D(n18383), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][28]~FF  (.D(n18382), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][29]~FF  (.D(n18381), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][30]~FF  (.D(n18380), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[25][31]~FF  (.D(n18379), .CE(ceg_net51309), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[25][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[25][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[25][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[25][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[25][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[25][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[25][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[25][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][8]~FF  (.D(n18435), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][9]~FF  (.D(n18434), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][10]~FF  (.D(n18433), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][11]~FF  (.D(n18432), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][12]~FF  (.D(n18431), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][13]~FF  (.D(n18430), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][14]~FF  (.D(n18429), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][15]~FF  (.D(n18428), .CE(ceg_net46504), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][16]~FF  (.D(n18427), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][17]~FF  (.D(n18426), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][18]~FF  (.D(n18425), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][19]~FF  (.D(n18424), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][20]~FF  (.D(n18423), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][21]~FF  (.D(n18422), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][22]~FF  (.D(n18421), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][23]~FF  (.D(n18420), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][24]~FF  (.D(n18419), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][25]~FF  (.D(n18418), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][26]~FF  (.D(n18417), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][27]~FF  (.D(n18416), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][28]~FF  (.D(n18415), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][29]~FF  (.D(n18414), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][30]~FF  (.D(n18413), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[26][31]~FF  (.D(n18412), .CE(ceg_net51373), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[26][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[26][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[26][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[26][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[26][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[26][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[26][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[26][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][8]~FF  (.D(n18468), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][9]~FF  (.D(n18467), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][10]~FF  (.D(n18466), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][11]~FF  (.D(n18465), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][12]~FF  (.D(n18464), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][13]~FF  (.D(n18463), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][14]~FF  (.D(n18462), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][15]~FF  (.D(n18461), .CE(ceg_net46696), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][16]~FF  (.D(n18460), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][17]~FF  (.D(n18459), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][18]~FF  (.D(n18458), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][19]~FF  (.D(n18457), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][20]~FF  (.D(n18456), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][21]~FF  (.D(n18455), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][22]~FF  (.D(n18454), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][23]~FF  (.D(n18453), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][24]~FF  (.D(n18452), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][25]~FF  (.D(n18451), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][26]~FF  (.D(n18450), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][27]~FF  (.D(n18449), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][28]~FF  (.D(n18448), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][29]~FF  (.D(n18447), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][30]~FF  (.D(n18446), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[27][31]~FF  (.D(n18445), .CE(ceg_net51437), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[27][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[27][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[27][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[27][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[27][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[27][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[27][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[27][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][8]~FF  (.D(n18501), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][9]~FF  (.D(n18500), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][10]~FF  (.D(n18499), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][11]~FF  (.D(n18498), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][12]~FF  (.D(n18497), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][13]~FF  (.D(n18496), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][14]~FF  (.D(n18495), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][15]~FF  (.D(n18494), .CE(ceg_net46888), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][16]~FF  (.D(n18493), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][17]~FF  (.D(n18492), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][18]~FF  (.D(n18491), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][19]~FF  (.D(n18490), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][20]~FF  (.D(n18489), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][21]~FF  (.D(n18488), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][22]~FF  (.D(n18487), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][23]~FF  (.D(n18486), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][24]~FF  (.D(n18485), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][25]~FF  (.D(n18484), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][26]~FF  (.D(n18483), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][27]~FF  (.D(n18482), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][28]~FF  (.D(n18481), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][29]~FF  (.D(n18480), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][30]~FF  (.D(n18479), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[28][31]~FF  (.D(n18478), .CE(ceg_net51501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[28][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[28][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[28][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[28][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[28][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[28][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[28][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[28][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][8]~FF  (.D(n18534), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][9]~FF  (.D(n18533), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][10]~FF  (.D(n18532), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][11]~FF  (.D(n18531), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][12]~FF  (.D(n18530), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][13]~FF  (.D(n18529), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][14]~FF  (.D(n18528), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][15]~FF  (.D(n18527), .CE(ceg_net47080), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][16]~FF  (.D(n18526), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][17]~FF  (.D(n18525), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][18]~FF  (.D(n18524), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][19]~FF  (.D(n18523), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][20]~FF  (.D(n18522), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][21]~FF  (.D(n18521), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][22]~FF  (.D(n18520), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][23]~FF  (.D(n18519), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][24]~FF  (.D(n18518), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][25]~FF  (.D(n18517), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][26]~FF  (.D(n18516), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][27]~FF  (.D(n18515), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][28]~FF  (.D(n18514), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][29]~FF  (.D(n18513), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][30]~FF  (.D(n18512), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[29][31]~FF  (.D(n18511), .CE(ceg_net51565), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[29][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[29][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[29][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[29][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[29][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[29][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[29][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[29][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][8]~FF  (.D(n18567), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][9]~FF  (.D(n18566), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][10]~FF  (.D(n18565), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][11]~FF  (.D(n18564), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][12]~FF  (.D(n18563), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][13]~FF  (.D(n18562), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][14]~FF  (.D(n18561), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][15]~FF  (.D(n18560), .CE(ceg_net47272), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][16]~FF  (.D(n18559), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][17]~FF  (.D(n18558), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][18]~FF  (.D(n18557), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][19]~FF  (.D(n18556), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][20]~FF  (.D(n18555), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][21]~FF  (.D(n18554), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][22]~FF  (.D(n18553), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][23]~FF  (.D(n18552), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][24]~FF  (.D(n18551), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][25]~FF  (.D(n18550), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][26]~FF  (.D(n18549), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][27]~FF  (.D(n18548), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][28]~FF  (.D(n18547), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][29]~FF  (.D(n18546), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][30]~FF  (.D(n18545), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[30][31]~FF  (.D(n18544), .CE(ceg_net51629), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[30][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[30][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[30][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[30][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[30][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[30][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[30][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[30][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][8]~FF  (.D(n18600), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][8]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][8]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][8]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][8]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][8]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][8]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][9]~FF  (.D(n18599), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][9]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][9]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][9]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][9]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][9]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][9]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][10]~FF  (.D(n18598), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][10]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][10]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][10]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][10]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][10]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][10]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][11]~FF  (.D(n18597), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][11]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][11]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][11]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][11]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][11]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][11]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][12]~FF  (.D(n18596), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][12]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][12]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][12]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][12]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][12]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][12]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][13]~FF  (.D(n18595), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][13]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][13]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][13]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][13]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][13]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][13]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][14]~FF  (.D(n18594), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][14]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][14]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][14]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][14]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][14]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][14]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][15]~FF  (.D(n18593), .CE(ceg_net47464), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][15]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][15]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][15]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][15]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][15]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][15]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][16]~FF  (.D(n18592), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][16]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][16]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][16]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][16]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][16]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][16]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][17]~FF  (.D(n18591), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][17]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][17]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][17]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][17]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][17]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][17]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][18]~FF  (.D(n18590), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][18]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][18]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][18]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][18]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][18]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][18]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][19]~FF  (.D(n18589), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][19]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][19]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][19]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][19]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][19]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][19]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][20]~FF  (.D(n18588), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][20]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][20]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][20]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][20]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][20]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][20]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][21]~FF  (.D(n18587), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][21]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][21]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][21]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][21]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][21]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][21]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][22]~FF  (.D(n18586), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][22]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][22]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][22]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][22]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][22]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][22]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][23]~FF  (.D(n18585), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][23]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][23]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][23]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][23]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][23]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][23]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][24]~FF  (.D(n18584), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][24]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][24]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][24]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][24]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][24]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][24]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][25]~FF  (.D(n18583), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][25]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][25]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][25]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][25]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][25]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][25]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][26]~FF  (.D(n18582), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][26]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][26]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][26]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][26]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][26]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][26]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][27]~FF  (.D(n18581), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][27]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][27]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][27]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][27]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][27]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][27]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][28]~FF  (.D(n18580), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][28]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][28]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][28]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][28]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][28]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][28]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][29]~FF  (.D(n18579), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][29]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][29]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][29]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][29]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][29]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][29]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][30]~FF  (.D(n18578), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][30]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][30]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][30]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][30]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][30]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][30]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XI[31][31]~FF  (.D(n18577), .CE(ceg_net51753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XI[31][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XI[31][31]~FF .CLK_POLARITY = 1'b1;
    defparam \XI[31][31]~FF .CE_POLARITY = 1'b1;
    defparam \XI[31][31]~FF .SR_POLARITY = 1'b1;
    defparam \XI[31][31]~FF .D_POLARITY = 1'b1;
    defparam \XI[31][31]~FF .SR_SYNC = 1'b1;
    defparam \XI[31][31]~FF .SR_VALUE = 1'b0;
    defparam \XI[31][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][1]~FF  (.D(n19663), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][2]~FF  (.D(n19662), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][3]~FF  (.D(n19661), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][4]~FF  (.D(n19660), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][5]~FF  (.D(n19659), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][6]~FF  (.D(n19658), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[0][7]~FF  (.D(n19657), .CE(ceg_net27233), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[0][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[0][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[0][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][1]~FF  (.D(n19663), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][2]~FF  (.D(n19662), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][3]~FF  (.D(n19661), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][4]~FF  (.D(n19660), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][5]~FF  (.D(n19659), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][6]~FF  (.D(n19658), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[1][7]~FF  (.D(n19657), .CE(ceg_net27485), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[1][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[1][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[1][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][1]~FF  (.D(n19663), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][2]~FF  (.D(n19662), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][3]~FF  (.D(n19661), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][4]~FF  (.D(n19660), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][5]~FF  (.D(n19659), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][6]~FF  (.D(n19658), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[2][7]~FF  (.D(n19657), .CE(ceg_net27737), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[2][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[2][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[2][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[2][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[2][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[2][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[2][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[2][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][1]~FF  (.D(n19663), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][2]~FF  (.D(n19662), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][3]~FF  (.D(n19661), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][4]~FF  (.D(n19660), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][5]~FF  (.D(n19659), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][6]~FF  (.D(n19658), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[3][7]~FF  (.D(n19657), .CE(ceg_net27989), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[3][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[3][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[3][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[3][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[3][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[3][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[3][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[3][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][1]~FF  (.D(n19663), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][2]~FF  (.D(n19662), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][3]~FF  (.D(n19661), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][4]~FF  (.D(n19660), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][5]~FF  (.D(n19659), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][6]~FF  (.D(n19658), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[4][7]~FF  (.D(n19657), .CE(ceg_net28241), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[4][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[4][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[4][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[4][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[4][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[4][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[4][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[4][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][1]~FF  (.D(n19663), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][2]~FF  (.D(n19662), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][3]~FF  (.D(n19661), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][4]~FF  (.D(n19660), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][5]~FF  (.D(n19659), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][6]~FF  (.D(n19658), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[5][7]~FF  (.D(n19657), .CE(ceg_net28493), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[5][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[5][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[5][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[5][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[5][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[5][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[5][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[5][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][1]~FF  (.D(n19663), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][2]~FF  (.D(n19662), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][3]~FF  (.D(n19661), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][4]~FF  (.D(n19660), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][5]~FF  (.D(n19659), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][6]~FF  (.D(n19658), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[6][7]~FF  (.D(n19657), .CE(ceg_net28745), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[6][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[6][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[6][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[6][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[6][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[6][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[6][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[6][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][1]~FF  (.D(n19663), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][2]~FF  (.D(n19662), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][3]~FF  (.D(n19661), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][4]~FF  (.D(n19660), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][5]~FF  (.D(n19659), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][6]~FF  (.D(n19658), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[7][7]~FF  (.D(n19657), .CE(ceg_net28997), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[7][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[7][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[7][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[7][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[7][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[7][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[7][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[7][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][1]~FF  (.D(n19663), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][2]~FF  (.D(n19662), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][3]~FF  (.D(n19661), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][4]~FF  (.D(n19660), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][5]~FF  (.D(n19659), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][6]~FF  (.D(n19658), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[8][7]~FF  (.D(n19657), .CE(ceg_net29249), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[8][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[8][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[8][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[8][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[8][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[8][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[8][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[8][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][1]~FF  (.D(n19663), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][2]~FF  (.D(n19662), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][3]~FF  (.D(n19661), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][4]~FF  (.D(n19660), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][5]~FF  (.D(n19659), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][6]~FF  (.D(n19658), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[9][7]~FF  (.D(n19657), .CE(ceg_net29501), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[9][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[9][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[9][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[9][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[9][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[9][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[9][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[9][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][1]~FF  (.D(n19663), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][2]~FF  (.D(n19662), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][3]~FF  (.D(n19661), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][4]~FF  (.D(n19660), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][5]~FF  (.D(n19659), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][6]~FF  (.D(n19658), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[10][7]~FF  (.D(n19657), .CE(ceg_net29753), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[10][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[10][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[10][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[10][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[10][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[10][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[10][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[10][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][1]~FF  (.D(n19663), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][2]~FF  (.D(n19662), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][3]~FF  (.D(n19661), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][4]~FF  (.D(n19660), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][5]~FF  (.D(n19659), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][6]~FF  (.D(n19658), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[11][7]~FF  (.D(n19657), .CE(ceg_net30005), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[11][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[11][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[11][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[11][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[11][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[11][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[11][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[11][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][1]~FF  (.D(n19663), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][2]~FF  (.D(n19662), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][3]~FF  (.D(n19661), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][4]~FF  (.D(n19660), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][5]~FF  (.D(n19659), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][6]~FF  (.D(n19658), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[12][7]~FF  (.D(n19657), .CE(ceg_net30257), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[12][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[12][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[12][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[12][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[12][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[12][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[12][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[12][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][1]~FF  (.D(n19663), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][2]~FF  (.D(n19662), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][3]~FF  (.D(n19661), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][4]~FF  (.D(n19660), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][5]~FF  (.D(n19659), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][6]~FF  (.D(n19658), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[13][7]~FF  (.D(n19657), .CE(ceg_net30509), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[13][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[13][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[13][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[13][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[13][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[13][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[13][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[13][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][1]~FF  (.D(n19663), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][2]~FF  (.D(n19662), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][3]~FF  (.D(n19661), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][4]~FF  (.D(n19660), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][5]~FF  (.D(n19659), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][6]~FF  (.D(n19658), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[14][7]~FF  (.D(n19657), .CE(ceg_net30761), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[14][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[14][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[14][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[14][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[14][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[14][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[14][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[14][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][1]~FF  (.D(n19663), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][2]~FF  (.D(n19662), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][3]~FF  (.D(n19661), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][4]~FF  (.D(n19660), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][5]~FF  (.D(n19659), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][6]~FF  (.D(n19658), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[15][7]~FF  (.D(n19657), .CE(ceg_net31013), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[15][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[15][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[15][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[15][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[15][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[15][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[15][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[15][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][1]~FF  (.D(n19663), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][2]~FF  (.D(n19662), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][3]~FF  (.D(n19661), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][4]~FF  (.D(n19660), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][5]~FF  (.D(n19659), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][6]~FF  (.D(n19658), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[16][7]~FF  (.D(n19657), .CE(ceg_net31265), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[16][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[16][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[16][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[16][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[16][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[16][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[16][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[16][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][1]~FF  (.D(n19663), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][2]~FF  (.D(n19662), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][3]~FF  (.D(n19661), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][4]~FF  (.D(n19660), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][5]~FF  (.D(n19659), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][6]~FF  (.D(n19658), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[17][7]~FF  (.D(n19657), .CE(ceg_net31517), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[17][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[17][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[17][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[17][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[17][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[17][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[17][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[17][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][1]~FF  (.D(n19663), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][2]~FF  (.D(n19662), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][3]~FF  (.D(n19661), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][4]~FF  (.D(n19660), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][5]~FF  (.D(n19659), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][6]~FF  (.D(n19658), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[18][7]~FF  (.D(n19657), .CE(ceg_net31769), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[18][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[18][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[18][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[18][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[18][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[18][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[18][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[18][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][1]~FF  (.D(n19663), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][2]~FF  (.D(n19662), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][3]~FF  (.D(n19661), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][4]~FF  (.D(n19660), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][5]~FF  (.D(n19659), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][6]~FF  (.D(n19658), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[19][7]~FF  (.D(n19657), .CE(ceg_net32021), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[19][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[19][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[19][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[19][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[19][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[19][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[19][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[19][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][1]~FF  (.D(n19663), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][2]~FF  (.D(n19662), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][3]~FF  (.D(n19661), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][4]~FF  (.D(n19660), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][5]~FF  (.D(n19659), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][6]~FF  (.D(n19658), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[20][7]~FF  (.D(n19657), .CE(ceg_net32273), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[20][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[20][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[20][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[20][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[20][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[20][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[20][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[20][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][1]~FF  (.D(n19663), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][2]~FF  (.D(n19662), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][3]~FF  (.D(n19661), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][4]~FF  (.D(n19660), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][5]~FF  (.D(n19659), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][6]~FF  (.D(n19658), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[21][7]~FF  (.D(n19657), .CE(ceg_net32525), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[21][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[21][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[21][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[21][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[21][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[21][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[21][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[21][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][1]~FF  (.D(n19663), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][2]~FF  (.D(n19662), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][3]~FF  (.D(n19661), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][4]~FF  (.D(n19660), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][5]~FF  (.D(n19659), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][6]~FF  (.D(n19658), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[22][7]~FF  (.D(n19657), .CE(ceg_net32777), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[22][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[22][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[22][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[22][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[22][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[22][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[22][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[22][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][1]~FF  (.D(n19663), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][2]~FF  (.D(n19662), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][3]~FF  (.D(n19661), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][4]~FF  (.D(n19660), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][5]~FF  (.D(n19659), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][6]~FF  (.D(n19658), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[23][7]~FF  (.D(n19657), .CE(ceg_net33029), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[23][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[23][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[23][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[23][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[23][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[23][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[23][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[23][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][1]~FF  (.D(n19663), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][2]~FF  (.D(n19662), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][3]~FF  (.D(n19661), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][4]~FF  (.D(n19660), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][5]~FF  (.D(n19659), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][6]~FF  (.D(n19658), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[24][7]~FF  (.D(n19657), .CE(ceg_net33281), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[24][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[24][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[24][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[24][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[24][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[24][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[24][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[24][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][1]~FF  (.D(n19663), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][2]~FF  (.D(n19662), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][3]~FF  (.D(n19661), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][4]~FF  (.D(n19660), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][5]~FF  (.D(n19659), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][6]~FF  (.D(n19658), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[25][7]~FF  (.D(n19657), .CE(ceg_net33533), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[25][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[25][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[25][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[25][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[25][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[25][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[25][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[25][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][1]~FF  (.D(n19663), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][2]~FF  (.D(n19662), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][3]~FF  (.D(n19661), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][4]~FF  (.D(n19660), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][5]~FF  (.D(n19659), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][6]~FF  (.D(n19658), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[26][7]~FF  (.D(n19657), .CE(ceg_net33785), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[26][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[26][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[26][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[26][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[26][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[26][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[26][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[26][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][1]~FF  (.D(n19663), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][2]~FF  (.D(n19662), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][3]~FF  (.D(n19661), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][4]~FF  (.D(n19660), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][5]~FF  (.D(n19659), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][6]~FF  (.D(n19658), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[27][7]~FF  (.D(n19657), .CE(ceg_net34037), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[27][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[27][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[27][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[27][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[27][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[27][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[27][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[27][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][1]~FF  (.D(n19663), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][2]~FF  (.D(n19662), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][3]~FF  (.D(n19661), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][4]~FF  (.D(n19660), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][5]~FF  (.D(n19659), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][6]~FF  (.D(n19658), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[28][7]~FF  (.D(n19657), .CE(ceg_net34289), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[28][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[28][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[28][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[28][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[28][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[28][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[28][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[28][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][1]~FF  (.D(n19663), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][2]~FF  (.D(n19662), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][3]~FF  (.D(n19661), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][4]~FF  (.D(n19660), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][5]~FF  (.D(n19659), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][6]~FF  (.D(n19658), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[29][7]~FF  (.D(n19657), .CE(ceg_net34541), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[29][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[29][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[29][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[29][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[29][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[29][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[29][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[29][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][1]~FF  (.D(n19663), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][2]~FF  (.D(n19662), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][3]~FF  (.D(n19661), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][4]~FF  (.D(n19660), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][5]~FF  (.D(n19659), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][6]~FF  (.D(n19658), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[30][7]~FF  (.D(n19657), .CE(ceg_net34793), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[30][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[30][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[30][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[30][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[30][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[30][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[30][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[30][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][1]~FF  (.D(n19663), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][1]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][1]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][1]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][1]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][1]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][1]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][2]~FF  (.D(n19662), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][2]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][2]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][2]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][2]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][2]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][2]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][3]~FF  (.D(n19661), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][3]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][3]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][3]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][3]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][3]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][3]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][4]~FF  (.D(n19660), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][4]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][4]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][4]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][4]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][4]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][4]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][5]~FF  (.D(n19659), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][5]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][5]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][5]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][5]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][5]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][5]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][6]~FF  (.D(n19658), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][6]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][6]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][6]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][6]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][6]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][6]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XII[31][7]~FF  (.D(n19657), .CE(ceg_net18979), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\XII[31][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(636)
    defparam \XII[31][7]~FF .CLK_POLARITY = 1'b1;
    defparam \XII[31][7]~FF .CE_POLARITY = 1'b1;
    defparam \XII[31][7]~FF .SR_POLARITY = 1'b1;
    defparam \XII[31][7]~FF .D_POLARITY = 1'b1;
    defparam \XII[31][7]~FF .SR_SYNC = 1'b1;
    defparam \XII[31][7]~FF .SR_VALUE = 1'b0;
    defparam \XII[31][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__4494 (.I0(STAGE2_EN), .I1(n51770), .O(n2954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4494.LUTMASK = 16'h8888;
    EFX_ADD \add_183/i1  (.I0(\ARG1[0] ), .I1(\ARG2[0] ), .CI(1'b0), .O(n8), 
            .CO(n9)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i1 .I0_POLARITY = 1'b1;
    defparam \add_183/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i1  (.I0(\ARG1[0] ), .I1(\ARG3[0] ), .CI(1'b0), .O(n32), 
            .CO(n33)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i1 .I0_POLARITY = 1'b1;
    defparam \add_207/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_184/add_2/i1  (.I0(\ARG1[0] ), .I1(\ARG2[0] ), .CI(n5921), 
            .O(n39), .CO(n40)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i32  (.I0(\ARG1[31] ), .I1(\ARG2[31] ), .CI(n5922), 
            .O(n1341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i32 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i31  (.I0(\ARG1[30] ), .I1(\ARG2[30] ), .CI(n5923), 
            .O(n1342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i31 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i30  (.I0(\ARG1[29] ), .I1(\ARG2[29] ), .CI(n5924), 
            .O(n1343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i30 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i29  (.I0(\ARG1[28] ), .I1(\ARG2[28] ), .CI(n5925), 
            .O(n1344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i29 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i28  (.I0(\ARG1[27] ), .I1(\ARG2[27] ), .CI(n5926), 
            .O(n1345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i27  (.I0(\ARG1[26] ), .I1(\ARG2[26] ), .CI(n5927), 
            .O(n1346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i26  (.I0(\ARG1[25] ), .I1(\ARG2[25] ), .CI(n5928), 
            .O(n1347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i25  (.I0(\ARG1[24] ), .I1(\ARG2[24] ), .CI(n5929), 
            .O(n1348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i24  (.I0(\ARG1[23] ), .I1(\ARG2[23] ), .CI(n5930), 
            .O(n1349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i23  (.I0(\ARG1[22] ), .I1(\ARG2[22] ), .CI(n5931), 
            .O(n1350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i22  (.I0(\ARG1[21] ), .I1(\ARG2[21] ), .CI(n5932), 
            .O(n1351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i21  (.I0(\ARG1[20] ), .I1(\ARG2[20] ), .CI(n5933), 
            .O(n1352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i20  (.I0(\ARG1[19] ), .I1(\ARG2[19] ), .CI(n5934), 
            .O(n1353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i19  (.I0(\ARG1[18] ), .I1(\ARG2[18] ), .CI(n5935), 
            .O(n1354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i18  (.I0(\ARG1[17] ), .I1(\ARG2[17] ), .CI(n5936), 
            .O(n1355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i17  (.I0(\ARG1[16] ), .I1(\ARG2[16] ), .CI(n5937), 
            .O(n1356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i16  (.I0(\ARG1[15] ), .I1(\ARG2[15] ), .CI(n5938), 
            .O(n1357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i15  (.I0(\ARG1[14] ), .I1(\ARG2[14] ), .CI(n5939), 
            .O(n1358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i14  (.I0(\ARG1[13] ), .I1(\ARG2[13] ), .CI(n5940), 
            .O(n1359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i13  (.I0(\ARG1[12] ), .I1(\ARG2[12] ), .CI(n5941), 
            .O(n1360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i12  (.I0(\ARG1[11] ), .I1(\ARG2[11] ), .CI(n5942), 
            .O(n1361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i11  (.I0(\ARG1[10] ), .I1(\ARG2[10] ), .CI(n5943), 
            .O(n1362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i10  (.I0(\ARG1[9] ), .I1(\ARG2[9] ), .CI(n5944), 
            .O(n1363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i9  (.I0(\ARG1[8] ), .I1(\ARG2[8] ), .CI(n5945), 
            .O(n1364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i8  (.I0(\ARG1[7] ), .I1(\ARG2[7] ), .CI(n5946), 
            .O(n1365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i7  (.I0(\ARG1[6] ), .I1(\ARG2[6] ), .CI(n5947), 
            .O(n1366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i6  (.I0(\ARG1[5] ), .I1(\ARG2[5] ), .CI(n5948), 
            .O(n1367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i5  (.I0(\ARG1[4] ), .I1(\ARG2[4] ), .CI(n5949), 
            .O(n1368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i4  (.I0(\ARG1[3] ), .I1(\ARG2[3] ), .CI(n5950), 
            .O(n1369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i3  (.I0(\ARG1[2] ), .I1(\ARG2[2] ), .CI(n5951), 
            .O(n1370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \sub_184/add_2/i2  (.I0(\ARG1[1] ), .I1(\ARG2[1] ), .CI(n40), 
            .O(n1371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \sub_184/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \sub_184/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \add_207/i10  (.I0(\ARG1[9] ), .I1(\ARG3[9] ), .CI(n1374), 
            .O(n1372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i10 .I0_POLARITY = 1'b1;
    defparam \add_207/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i9  (.I0(\ARG1[8] ), .I1(\ARG3[8] ), .CI(n1376), 
            .O(n1373), .CO(n1374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i9 .I0_POLARITY = 1'b1;
    defparam \add_207/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i8  (.I0(\ARG1[7] ), .I1(\ARG3[7] ), .CI(n1378), 
            .O(n1375), .CO(n1376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i8 .I0_POLARITY = 1'b1;
    defparam \add_207/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i7  (.I0(\ARG1[6] ), .I1(\ARG3[6] ), .CI(n1380), 
            .O(n1377), .CO(n1378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i7 .I0_POLARITY = 1'b1;
    defparam \add_207/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i6  (.I0(\ARG1[5] ), .I1(\ARG3[5] ), .CI(n1382), 
            .O(n1379), .CO(n1380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i6 .I0_POLARITY = 1'b1;
    defparam \add_207/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i5  (.I0(\ARG1[4] ), .I1(\ARG3[4] ), .CI(n1384), 
            .O(n1381), .CO(n1382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i5 .I0_POLARITY = 1'b1;
    defparam \add_207/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i4  (.I0(\ARG1[3] ), .I1(\ARG3[3] ), .CI(n1386), 
            .O(n1383), .CO(n1384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i4 .I0_POLARITY = 1'b1;
    defparam \add_207/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i3  (.I0(\ARG1[2] ), .I1(\ARG3[2] ), .CI(n1388), 
            .O(n1385), .CO(n1386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i3 .I0_POLARITY = 1'b1;
    defparam \add_207/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_207/i2  (.I0(\ARG1[1] ), .I1(\ARG3[1] ), .CI(n33), .O(n1387), 
            .CO(n1388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(583)
    defparam \add_207/i2 .I0_POLARITY = 1'b1;
    defparam \add_207/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i32  (.I0(\ARG1[31] ), .I1(\ARG2[31] ), .CI(n1391), 
            .O(n1389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i32 .I0_POLARITY = 1'b1;
    defparam \add_183/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i31  (.I0(\ARG1[30] ), .I1(\ARG2[30] ), .CI(n1393), 
            .O(n1390), .CO(n1391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i31 .I0_POLARITY = 1'b1;
    defparam \add_183/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i30  (.I0(\ARG1[29] ), .I1(\ARG2[29] ), .CI(n1395), 
            .O(n1392), .CO(n1393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i30 .I0_POLARITY = 1'b1;
    defparam \add_183/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i29  (.I0(\ARG1[28] ), .I1(\ARG2[28] ), .CI(n1397), 
            .O(n1394), .CO(n1395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i29 .I0_POLARITY = 1'b1;
    defparam \add_183/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i28  (.I0(\ARG1[27] ), .I1(\ARG2[27] ), .CI(n1399), 
            .O(n1396), .CO(n1397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i28 .I0_POLARITY = 1'b1;
    defparam \add_183/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i27  (.I0(\ARG1[26] ), .I1(\ARG2[26] ), .CI(n1401), 
            .O(n1398), .CO(n1399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i27 .I0_POLARITY = 1'b1;
    defparam \add_183/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i26  (.I0(\ARG1[25] ), .I1(\ARG2[25] ), .CI(n1403), 
            .O(n1400), .CO(n1401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i26 .I0_POLARITY = 1'b1;
    defparam \add_183/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i25  (.I0(\ARG1[24] ), .I1(\ARG2[24] ), .CI(n1405), 
            .O(n1402), .CO(n1403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i25 .I0_POLARITY = 1'b1;
    defparam \add_183/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i24  (.I0(\ARG1[23] ), .I1(\ARG2[23] ), .CI(n1407), 
            .O(n1404), .CO(n1405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i24 .I0_POLARITY = 1'b1;
    defparam \add_183/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i23  (.I0(\ARG1[22] ), .I1(\ARG2[22] ), .CI(n1409), 
            .O(n1406), .CO(n1407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i23 .I0_POLARITY = 1'b1;
    defparam \add_183/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i22  (.I0(\ARG1[21] ), .I1(\ARG2[21] ), .CI(n1411), 
            .O(n1408), .CO(n1409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i22 .I0_POLARITY = 1'b1;
    defparam \add_183/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i21  (.I0(\ARG1[20] ), .I1(\ARG2[20] ), .CI(n1413), 
            .O(n1410), .CO(n1411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i21 .I0_POLARITY = 1'b1;
    defparam \add_183/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i20  (.I0(\ARG1[19] ), .I1(\ARG2[19] ), .CI(n1415), 
            .O(n1412), .CO(n1413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i20 .I0_POLARITY = 1'b1;
    defparam \add_183/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i19  (.I0(\ARG1[18] ), .I1(\ARG2[18] ), .CI(n1417), 
            .O(n1414), .CO(n1415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i19 .I0_POLARITY = 1'b1;
    defparam \add_183/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i18  (.I0(\ARG1[17] ), .I1(\ARG2[17] ), .CI(n1419), 
            .O(n1416), .CO(n1417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i18 .I0_POLARITY = 1'b1;
    defparam \add_183/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i17  (.I0(\ARG1[16] ), .I1(\ARG2[16] ), .CI(n1421), 
            .O(n1418), .CO(n1419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i17 .I0_POLARITY = 1'b1;
    defparam \add_183/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i16  (.I0(\ARG1[15] ), .I1(\ARG2[15] ), .CI(n1423), 
            .O(n1420), .CO(n1421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i16 .I0_POLARITY = 1'b1;
    defparam \add_183/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i15  (.I0(\ARG1[14] ), .I1(\ARG2[14] ), .CI(n1425), 
            .O(n1422), .CO(n1423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i15 .I0_POLARITY = 1'b1;
    defparam \add_183/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i14  (.I0(\ARG1[13] ), .I1(\ARG2[13] ), .CI(n1427), 
            .O(n1424), .CO(n1425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i14 .I0_POLARITY = 1'b1;
    defparam \add_183/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i13  (.I0(\ARG1[12] ), .I1(\ARG2[12] ), .CI(n1429), 
            .O(n1426), .CO(n1427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i13 .I0_POLARITY = 1'b1;
    defparam \add_183/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i12  (.I0(\ARG1[11] ), .I1(\ARG2[11] ), .CI(n1431), 
            .O(n1428), .CO(n1429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i12 .I0_POLARITY = 1'b1;
    defparam \add_183/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i11  (.I0(\ARG1[10] ), .I1(\ARG2[10] ), .CI(n1433), 
            .O(n1430), .CO(n1431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i11 .I0_POLARITY = 1'b1;
    defparam \add_183/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i10  (.I0(\ARG1[9] ), .I1(\ARG2[9] ), .CI(n1435), 
            .O(n1432), .CO(n1433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i10 .I0_POLARITY = 1'b1;
    defparam \add_183/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i9  (.I0(\ARG1[8] ), .I1(\ARG2[8] ), .CI(n1437), 
            .O(n1434), .CO(n1435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i9 .I0_POLARITY = 1'b1;
    defparam \add_183/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i8  (.I0(\ARG1[7] ), .I1(\ARG2[7] ), .CI(n1439), 
            .O(n1436), .CO(n1437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i8 .I0_POLARITY = 1'b1;
    defparam \add_183/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i7  (.I0(\ARG1[6] ), .I1(\ARG2[6] ), .CI(n1441), 
            .O(n1438), .CO(n1439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i7 .I0_POLARITY = 1'b1;
    defparam \add_183/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i6  (.I0(\ARG1[5] ), .I1(\ARG2[5] ), .CI(n1443), 
            .O(n1440), .CO(n1441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i6 .I0_POLARITY = 1'b1;
    defparam \add_183/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i5  (.I0(\ARG1[4] ), .I1(\ARG2[4] ), .CI(n1445), 
            .O(n1442), .CO(n1443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i5 .I0_POLARITY = 1'b1;
    defparam \add_183/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i4  (.I0(\ARG1[3] ), .I1(\ARG2[3] ), .CI(n1447), 
            .O(n1444), .CO(n1445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i4 .I0_POLARITY = 1'b1;
    defparam \add_183/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i3  (.I0(\ARG1[2] ), .I1(\ARG2[2] ), .CI(n1449), 
            .O(n1446), .CO(n1447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i3 .I0_POLARITY = 1'b1;
    defparam \add_183/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_183/i2  (.I0(\ARG1[1] ), .I1(\ARG2[1] ), .CI(n9), .O(n1448), 
            .CO(n1449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(569)
    defparam \add_183/i2 .I0_POLARITY = 1'b1;
    defparam \add_183/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i32  (.I0(\PC[31] ), .I1(1'b0), .CI(n1452), .O(n1450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i32 .I0_POLARITY = 1'b1;
    defparam \add_24/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i31  (.I0(\PC[30] ), .I1(1'b0), .CI(n1454), .O(n1451), 
            .CO(n1452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i31 .I0_POLARITY = 1'b1;
    defparam \add_24/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i30  (.I0(\PC[29] ), .I1(1'b0), .CI(n1456), .O(n1453), 
            .CO(n1454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i30 .I0_POLARITY = 1'b1;
    defparam \add_24/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i29  (.I0(\PC[28] ), .I1(1'b0), .CI(n1458), .O(n1455), 
            .CO(n1456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i29 .I0_POLARITY = 1'b1;
    defparam \add_24/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i28  (.I0(\PC[27] ), .I1(1'b0), .CI(n1460), .O(n1457), 
            .CO(n1458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i28 .I0_POLARITY = 1'b1;
    defparam \add_24/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i27  (.I0(\PC[26] ), .I1(1'b0), .CI(n1462), .O(n1459), 
            .CO(n1460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i27 .I0_POLARITY = 1'b1;
    defparam \add_24/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i26  (.I0(\PC[25] ), .I1(1'b0), .CI(n1464), .O(n1461), 
            .CO(n1462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i26 .I0_POLARITY = 1'b1;
    defparam \add_24/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i25  (.I0(\PC[24] ), .I1(1'b0), .CI(n1466), .O(n1463), 
            .CO(n1464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i25 .I0_POLARITY = 1'b1;
    defparam \add_24/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i24  (.I0(\PC[23] ), .I1(1'b0), .CI(n1468), .O(n1465), 
            .CO(n1466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i24 .I0_POLARITY = 1'b1;
    defparam \add_24/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i23  (.I0(\PC[22] ), .I1(1'b0), .CI(n1470), .O(n1467), 
            .CO(n1468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i23 .I0_POLARITY = 1'b1;
    defparam \add_24/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i22  (.I0(\PC[21] ), .I1(1'b0), .CI(n1472), .O(n1469), 
            .CO(n1470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i22 .I0_POLARITY = 1'b1;
    defparam \add_24/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i21  (.I0(\PC[20] ), .I1(1'b0), .CI(n1474), .O(n1471), 
            .CO(n1472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i21 .I0_POLARITY = 1'b1;
    defparam \add_24/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i20  (.I0(\PC[19] ), .I1(1'b0), .CI(n1476), .O(n1473), 
            .CO(n1474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i20 .I0_POLARITY = 1'b1;
    defparam \add_24/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i19  (.I0(\PC[18] ), .I1(1'b0), .CI(n1478), .O(n1475), 
            .CO(n1476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i19 .I0_POLARITY = 1'b1;
    defparam \add_24/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i18  (.I0(\PC[17] ), .I1(1'b0), .CI(n1480), .O(n1477), 
            .CO(n1478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i18 .I0_POLARITY = 1'b1;
    defparam \add_24/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i17  (.I0(\PC[16] ), .I1(1'b0), .CI(n1482), .O(n1479), 
            .CO(n1480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i17 .I0_POLARITY = 1'b1;
    defparam \add_24/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i16  (.I0(\PC[15] ), .I1(1'b0), .CI(n1484), .O(n1481), 
            .CO(n1482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i16 .I0_POLARITY = 1'b1;
    defparam \add_24/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i15  (.I0(\PC[14] ), .I1(1'b0), .CI(n1486), .O(n1483), 
            .CO(n1484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i15 .I0_POLARITY = 1'b1;
    defparam \add_24/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i14  (.I0(\PC[13] ), .I1(1'b0), .CI(n1488), .O(n1485), 
            .CO(n1486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i14 .I0_POLARITY = 1'b1;
    defparam \add_24/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i13  (.I0(\PC[12] ), .I1(1'b0), .CI(n1490), .O(n1487), 
            .CO(n1488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i13 .I0_POLARITY = 1'b1;
    defparam \add_24/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i12  (.I0(\PC[11] ), .I1(1'b0), .CI(n1492), .O(n1489), 
            .CO(n1490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i12 .I0_POLARITY = 1'b1;
    defparam \add_24/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i11  (.I0(\PC[10] ), .I1(1'b0), .CI(n1494), .O(n1491), 
            .CO(n1492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i11 .I0_POLARITY = 1'b1;
    defparam \add_24/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i10  (.I0(\PC[9] ), .I1(1'b0), .CI(n1496), .O(n1493), 
            .CO(n1494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i10 .I0_POLARITY = 1'b1;
    defparam \add_24/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i9  (.I0(\PC[8] ), .I1(1'b0), .CI(n1498), .O(n1495), 
            .CO(n1496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i9 .I0_POLARITY = 1'b1;
    defparam \add_24/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i8  (.I0(\PC[7] ), .I1(1'b0), .CI(n1500), .O(n1497), 
            .CO(n1498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i8 .I0_POLARITY = 1'b1;
    defparam \add_24/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i7  (.I0(\PC[6] ), .I1(1'b0), .CI(n1502), .O(n1499), 
            .CO(n1500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i7 .I0_POLARITY = 1'b1;
    defparam \add_24/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i6  (.I0(\PC[5] ), .I1(1'b0), .CI(n1504), .O(n1501), 
            .CO(n1502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i6 .I0_POLARITY = 1'b1;
    defparam \add_24/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i5  (.I0(\PC[4] ), .I1(1'b0), .CI(n1506), .O(n1503), 
            .CO(n1504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i5 .I0_POLARITY = 1'b1;
    defparam \add_24/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i4  (.I0(\PC[3] ), .I1(1'b0), .CI(n1508), .O(n1505), 
            .CO(n1506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i4 .I0_POLARITY = 1'b1;
    defparam \add_24/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i3  (.I0(\PC[2] ), .I1(1'b0), .CI(n1510), .O(n1507), 
            .CO(n1508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i3 .I0_POLARITY = 1'b1;
    defparam \add_24/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_24/i2  (.I0(\PC[1] ), .I1(\PC[0] ), .CI(1'b0), .O(n1509), 
            .CO(n1510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // ../vhdl_packages/vhdl_2008/src/numeric_std-body.vhdl(496)
    defparam \add_24/i2 .I0_POLARITY = 1'b1;
    defparam \add_24/i2 .I1_POLARITY = 1'b0;
    EFX_RAM_5K USER_MEM__D$12 (.WCLK(\CLK~O ), .RCLK(\CLK~O ), .WCLKE(n30807), 
            .WE(MEM_STORE), .RE(n50476), .WDATA({\SAVE_DATA[7] , \SAVE_DATA[6] , 
            \SAVE_DATA[5] , \SAVE_DATA[4] }), .WADDR({\SAVE_ADDRESS[9] , 
            \SAVE_ADDRESS[8] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[5] , 
            \SAVE_ADDRESS[4] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[1] , 
            \SAVE_ADDRESS[0] }), .RADDR({n1432, n1434, n1436, n1438, 
            n1440, n1442, n1444, n1446, n1448, n8}), .RDATA({\LOAD_DATA[7] , 
            \LOAD_DATA[6] , \LOAD_DATA[5] , \LOAD_DATA[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b0, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(234)
    defparam USER_MEM__D$12.READ_WIDTH = 4;
    defparam USER_MEM__D$12.WRITE_WIDTH = 4;
    defparam USER_MEM__D$12.WCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$12.WCLKE_POLARITY = 1'b1;
    defparam USER_MEM__D$12.WE_POLARITY = 1'b1;
    defparam USER_MEM__D$12.RCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$12.RE_POLARITY = 1'b0;
    defparam USER_MEM__D$12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$12.OUTPUT_REG = 1'b0;
    defparam USER_MEM__D$12.WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K PROG_MEM__D$b12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51830, 
            n51834})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h840820A50848840840030819405230819520000000003000000000000207BA3E, INIT_1=256'h0000000860B68840B64A61860840861010400000040404800000000000070A40, INIT_2=256'h0000000000400000000000021000000000000000000000800840000800040840, INIT_3=256'h2A4921030C0C00800202150010000000010200210212258310A1021260000048, INIT_4=256'h08430210C12101480C0010001010944004800814448040040B040518718D0400, INIT_5=256'h40200000C40C48A40C5A842A50C4084202841040004162009BA8841000006816, INIT_6=256'h92400A0280F8772B02880404408000484002406C840020100102480402CC4C4A, INIT_7=256'h0804000000000000000000048204068100891220840841990B0024024301D111, INIT_8=256'h840820A50848840840030819405230819520000000003000000000000207BA3E, INIT_9=256'h0000000860B68840B64A61860840861010400000040404800000000000070A40, INIT_A=256'h0000000000400000000000021000000000000000000000800840000800040840, INIT_B=256'h2A4921030C0C00800202150010000000010200210212258310A1021260000048, INIT_C=256'h08430210C12101480C0010001010944004800814448040040B040518718D0400, INIT_D=256'h40200000C40C48A40C5A842A50C4084202841040004162009BA8841000006816, INIT_E=256'h92400A0280F8772B02880404408000484002406C840020100102480402CC4C4A, INIT_F=256'h0804000000000000000000048204068100891220840841990B0024024301D111, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$b12.READ_WIDTH = 2;
    defparam PROG_MEM__D$b12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$b12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$b12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$b12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$b12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$b12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$b12.INIT_0 = 256'h840820A50848840840030819405230819520000000003000000000000207BA3E;
    defparam PROG_MEM__D$b12.INIT_1 = 256'h0000000860B68840B64A61860840861010400000040404800000000000070A40;
    defparam PROG_MEM__D$b12.INIT_2 = 256'h0000000000400000000000021000000000000000000000800840000800040840;
    defparam PROG_MEM__D$b12.INIT_3 = 256'h2A4921030C0C00800202150010000000010200210212258310A1021260000048;
    defparam PROG_MEM__D$b12.INIT_4 = 256'h08430210C12101480C0010001010944004800814448040040B040518718D0400;
    defparam PROG_MEM__D$b12.INIT_5 = 256'h40200000C40C48A40C5A842A50C4084202841040004162009BA8841000006816;
    defparam PROG_MEM__D$b12.INIT_6 = 256'h92400A0280F8772B02880404408000484002406C840020100102480402CC4C4A;
    defparam PROG_MEM__D$b12.INIT_7 = 256'h0804000000000000000000048204068100891220840841990B0024024301D111;
    defparam PROG_MEM__D$b12.INIT_8 = 256'h840820A50848840840030819405230819520000000003000000000000207BA3E;
    defparam PROG_MEM__D$b12.INIT_9 = 256'h0000000860B68840B64A61860840861010400000040404800000000000070A40;
    defparam PROG_MEM__D$b12.INIT_A = 256'h0000000000400000000000021000000000000000000000800840000800040840;
    defparam PROG_MEM__D$b12.INIT_B = 256'h2A4921030C0C00800202150010000000010200210212258310A1021260000048;
    defparam PROG_MEM__D$b12.INIT_C = 256'h08430210C12101480C0010001010944004800814448040040B040518718D0400;
    defparam PROG_MEM__D$b12.INIT_D = 256'h40200000C40C48A40C5A842A50C4084202841040004162009BA8841000006816;
    defparam PROG_MEM__D$b12.INIT_E = 256'h92400A0280F8772B02880404408000484002406C840020100102480402CC4C4A;
    defparam PROG_MEM__D$b12.INIT_F = 256'h0804000000000000000000048204068100891220840841990B0024024301D111;
    defparam PROG_MEM__D$b12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$b12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$b12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$b12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$b12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$b12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K USER_MEM__D$2 (.WCLK(\CLK~O ), .RCLK(\CLK~O ), .WCLKE(n30807), 
            .WE(MEM_STORE), .RE(n50476), .WDATA({\SAVE_DATA[3] , \SAVE_DATA[2] , 
            \SAVE_DATA[1] , \SAVE_DATA[0] }), .WADDR({\SAVE_ADDRESS[9] , 
            \SAVE_ADDRESS[8] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[5] , 
            \SAVE_ADDRESS[4] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[1] , 
            \SAVE_ADDRESS[0] }), .RADDR({n1432, n1434, n1436, n1438, 
            n1440, n1442, n1444, n1446, n1448, n8}), .RDATA({\LOAD_DATA[3] , 
            \LOAD_DATA[2] , \LOAD_DATA[1] , \LOAD_DATA[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b0, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(234)
    defparam USER_MEM__D$2.READ_WIDTH = 4;
    defparam USER_MEM__D$2.WRITE_WIDTH = 4;
    defparam USER_MEM__D$2.WCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$2.WCLKE_POLARITY = 1'b1;
    defparam USER_MEM__D$2.WE_POLARITY = 1'b1;
    defparam USER_MEM__D$2.RCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$2.RE_POLARITY = 1'b0;
    defparam USER_MEM__D$2.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$2.OUTPUT_REG = 1'b0;
    defparam USER_MEM__D$2.WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K PROG_MEM__D$o1 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51726, 
            n51730})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h18418618608419418603AA81965511A8181000000000C0000000000001511545, INIT_1=256'h00008003861A4184306186134184386000000000200800000000A00000186184, INIT_2=256'h0000000001000000000000040000020000000000000000000000000000000100, INIT_3=256'h1841020000200000000000140001021006106106106906106506106580000100, INIT_4=256'h40A01560A64940A4082004000000100C09D204000011000A600C1A01361221A4, INIT_5=256'h084000001841E4CCC0A40C4FC428428400080002480000000080080800018608, INIT_6=256'h830601008401800032000001008C4C000001540000C0003400503000040102D8, INIT_7=256'h00300000800002000008000081080080001020901A40124828280A408203C005, INIT_8=256'h18418618608419418603AA81965511A8181000000000C0000000000001511545, INIT_9=256'h00008003861A4184306186134184386000000000200800000000A00000186184, INIT_A=256'h0000000001000000000000040000020000000000000000000000000000000100, INIT_B=256'h1841020000200000000000140001021006106106106906106506106580000100, INIT_C=256'h40A01560A64940A4082004000000100C09D204000011000A600C1A01361221A4, INIT_D=256'h084000001841E4CCC0A40C4FC428428400080002480000000080080800018608, INIT_E=256'h830601008401800032000001008C4C000001540000C0003400503000040102D8, INIT_F=256'h00300000800002000008000081080080001020901A40124828280A408203C005, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$o1.READ_WIDTH = 2;
    defparam PROG_MEM__D$o1.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$o1.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$o1.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$o1.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$o1.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$o1.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$o1.INIT_0 = 256'h18418618608419418603AA81965511A8181000000000C0000000000001511545;
    defparam PROG_MEM__D$o1.INIT_1 = 256'h00008003861A4184306186134184386000000000200800000000A00000186184;
    defparam PROG_MEM__D$o1.INIT_2 = 256'h0000000001000000000000040000020000000000000000000000000000000100;
    defparam PROG_MEM__D$o1.INIT_3 = 256'h1841020000200000000000140001021006106106106906106506106580000100;
    defparam PROG_MEM__D$o1.INIT_4 = 256'h40A01560A64940A4082004000000100C09D204000011000A600C1A01361221A4;
    defparam PROG_MEM__D$o1.INIT_5 = 256'h084000001841E4CCC0A40C4FC428428400080002480000000080080800018608;
    defparam PROG_MEM__D$o1.INIT_6 = 256'h830601008401800032000001008C4C000001540000C0003400503000040102D8;
    defparam PROG_MEM__D$o1.INIT_7 = 256'h00300000800002000008000081080080001020901A40124828280A408203C005;
    defparam PROG_MEM__D$o1.INIT_8 = 256'h18418618608419418603AA81965511A8181000000000C0000000000001511545;
    defparam PROG_MEM__D$o1.INIT_9 = 256'h00008003861A4184306186134184386000000000200800000000A00000186184;
    defparam PROG_MEM__D$o1.INIT_A = 256'h0000000001000000000000040000020000000000000000000000000000000100;
    defparam PROG_MEM__D$o1.INIT_B = 256'h1841020000200000000000140001021006106106106906106506106580000100;
    defparam PROG_MEM__D$o1.INIT_C = 256'h40A01560A64940A4082004000000100C09D204000011000A600C1A01361221A4;
    defparam PROG_MEM__D$o1.INIT_D = 256'h084000001841E4CCC0A40C4FC428428400080002480000000080080800018608;
    defparam PROG_MEM__D$o1.INIT_E = 256'h830601008401800032000001008C4C000001540000C0003400503000040102D8;
    defparam PROG_MEM__D$o1.INIT_F = 256'h00300000800002000008000081080080001020901A40124828280A408203C005;
    defparam PROG_MEM__D$o1.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$o1.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$o1.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$o1.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$o1.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$o1.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K USER_MEM__D$c12 (.WCLK(\CLK~O ), .RCLK(\CLK~O ), .WCLKE(n30807), 
            .WE(MEM_STORE), .RE(n50476), .WDATA({\SAVE_DATA[16] , \SAVE_DATA[15] , 
            \SAVE_DATA[14] , \SAVE_DATA[13] , \SAVE_DATA[12] }), .WADDR({\SAVE_ADDRESS[9] , 
            \SAVE_ADDRESS[8] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[5] , 
            \SAVE_ADDRESS[4] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[1] , 
            \SAVE_ADDRESS[0] }), .RADDR({n1432, n1434, n1436, n1438, 
            n1440, n1442, n1444, n1446, n1448, n8}), .RDATA({\LOAD_DATA[16] , 
            \LOAD_DATA[15] , \LOAD_DATA[14] , \LOAD_DATA[13] , \LOAD_DATA[12] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b0, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(234)
    defparam USER_MEM__D$c12.READ_WIDTH = 5;
    defparam USER_MEM__D$c12.WRITE_WIDTH = 5;
    defparam USER_MEM__D$c12.WCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$c12.WCLKE_POLARITY = 1'b1;
    defparam USER_MEM__D$c12.WE_POLARITY = 1'b1;
    defparam USER_MEM__D$c12.RCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$c12.RE_POLARITY = 1'b0;
    defparam USER_MEM__D$c12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$c12.OUTPUT_REG = 1'b0;
    defparam USER_MEM__D$c12.WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K USER_MEM__D$d12 (.WCLK(\CLK~O ), .RCLK(\CLK~O ), .WCLKE(n30807), 
            .WE(MEM_STORE), .RE(n50476), .WDATA({\SAVE_DATA[21] , \SAVE_DATA[20] , 
            \SAVE_DATA[19] , \SAVE_DATA[18] , \SAVE_DATA[17] }), .WADDR({\SAVE_ADDRESS[9] , 
            \SAVE_ADDRESS[8] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[5] , 
            \SAVE_ADDRESS[4] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[1] , 
            \SAVE_ADDRESS[0] }), .RADDR({n1432, n1434, n1436, n1438, 
            n1440, n1442, n1444, n1446, n1448, n8}), .RDATA({\LOAD_DATA[21] , 
            \LOAD_DATA[20] , \LOAD_DATA[19] , \LOAD_DATA[18] , \LOAD_DATA[17] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b0, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(234)
    defparam USER_MEM__D$d12.READ_WIDTH = 5;
    defparam USER_MEM__D$d12.WRITE_WIDTH = 5;
    defparam USER_MEM__D$d12.WCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$d12.WCLKE_POLARITY = 1'b1;
    defparam USER_MEM__D$d12.WE_POLARITY = 1'b1;
    defparam USER_MEM__D$d12.RCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$d12.RE_POLARITY = 1'b0;
    defparam USER_MEM__D$d12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$d12.OUTPUT_REG = 1'b0;
    defparam USER_MEM__D$d12.WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K USER_MEM__D$e12 (.WCLK(\CLK~O ), .RCLK(\CLK~O ), .WCLKE(n30807), 
            .WE(MEM_STORE), .RE(n50476), .WDATA({\SAVE_DATA[26] , \SAVE_DATA[25] , 
            \SAVE_DATA[24] , \SAVE_DATA[23] , \SAVE_DATA[22] }), .WADDR({\SAVE_ADDRESS[9] , 
            \SAVE_ADDRESS[8] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[5] , 
            \SAVE_ADDRESS[4] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[1] , 
            \SAVE_ADDRESS[0] }), .RADDR({n1432, n1434, n1436, n1438, 
            n1440, n1442, n1444, n1446, n1448, n8}), .RDATA({\LOAD_DATA[26] , 
            \LOAD_DATA[25] , \LOAD_DATA[24] , \LOAD_DATA[23] , \LOAD_DATA[22] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b0, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(234)
    defparam USER_MEM__D$e12.READ_WIDTH = 5;
    defparam USER_MEM__D$e12.WRITE_WIDTH = 5;
    defparam USER_MEM__D$e12.WCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$e12.WCLKE_POLARITY = 1'b1;
    defparam USER_MEM__D$e12.WE_POLARITY = 1'b1;
    defparam USER_MEM__D$e12.RCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$e12.RE_POLARITY = 1'b0;
    defparam USER_MEM__D$e12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$e12.OUTPUT_REG = 1'b0;
    defparam USER_MEM__D$e12.WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K USER_MEM__D$f1 (.WCLK(\CLK~O ), .RCLK(\CLK~O ), .WCLKE(n30807), 
            .WE(MEM_STORE), .RE(n50476), .WDATA({\SAVE_DATA[31] , \SAVE_DATA[30] , 
            \SAVE_DATA[29] , \SAVE_DATA[28] , \SAVE_DATA[27] }), .WADDR({\SAVE_ADDRESS[9] , 
            \SAVE_ADDRESS[8] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[5] , 
            \SAVE_ADDRESS[4] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[1] , 
            \SAVE_ADDRESS[0] }), .RADDR({n1432, n1434, n1436, n1438, 
            n1440, n1442, n1444, n1446, n1448, n8}), .RDATA({\LOAD_DATA[31] , 
            \LOAD_DATA[30] , \LOAD_DATA[29] , \LOAD_DATA[28] , \LOAD_DATA[27] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b0, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(234)
    defparam USER_MEM__D$f1.READ_WIDTH = 5;
    defparam USER_MEM__D$f1.WRITE_WIDTH = 5;
    defparam USER_MEM__D$f1.WCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$f1.WCLKE_POLARITY = 1'b1;
    defparam USER_MEM__D$f1.WE_POLARITY = 1'b1;
    defparam USER_MEM__D$f1.RCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$f1.RE_POLARITY = 1'b0;
    defparam USER_MEM__D$f1.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$f1.OUTPUT_REG = 1'b0;
    defparam USER_MEM__D$f1.WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K PROG_MEM__D$n12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51734, 
            n51738})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h420051021020020001002EA0219544EA041000000000D000000000000D0AD8BB, INIT_1=256'h0000000021820040051001C40020461000000000000001004000000400021000, INIT_2=256'h0002102000100000000000000000000000040000000000001000040000000000, INIT_3=256'h0204010000100000008000200000102000844841940AC084A8408C2840010030, INIT_4=256'h0010821060000000205020832000022801010000000000001640050001421000, INIT_5=256'h300010004002800B402818C3B0420430010018400010011000404000000C6080, INIT_6=256'hC30A0232002B400C00D000003301B400818C38002013402001A020800B0030AC, INIT_7=256'h0401100100180400601001820025010200845400C504615056A040012103100B, INIT_8=256'h420051021020020001002EA0219544EA041000000000D000000000000D0AD8BB, INIT_9=256'h0000000021820040051001C40020461000000000000001004000000400021000, INIT_A=256'h0002102000100000000000000000000000040000000000001000040000000000, INIT_B=256'h0204010000100000008000200000102000844841940AC084A8408C2840010030, INIT_C=256'h0010821060000000205020832000022801010000000000001640050001421000, INIT_D=256'h300010004002800B402818C3B0420430010018400010011000404000000C6080, INIT_E=256'hC30A0232002B400C00D000003301B400818C38002013402001A020800B0030AC, INIT_F=256'h0401100100180400601001820025010200845400C504615056A040012103100B, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$n12.READ_WIDTH = 2;
    defparam PROG_MEM__D$n12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$n12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$n12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$n12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$n12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$n12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$n12.INIT_0 = 256'h420051021020020001002EA0219544EA041000000000D000000000000D0AD8BB;
    defparam PROG_MEM__D$n12.INIT_1 = 256'h0000000021820040051001C40020461000000000000001004000000400021000;
    defparam PROG_MEM__D$n12.INIT_2 = 256'h0002102000100000000000000000000000040000000000001000040000000000;
    defparam PROG_MEM__D$n12.INIT_3 = 256'h0204010000100000008000200000102000844841940AC084A8408C2840010030;
    defparam PROG_MEM__D$n12.INIT_4 = 256'h0010821060000000205020832000022801010000000000001640050001421000;
    defparam PROG_MEM__D$n12.INIT_5 = 256'h300010004002800B402818C3B0420430010018400010011000404000000C6080;
    defparam PROG_MEM__D$n12.INIT_6 = 256'hC30A0232002B400C00D000003301B400818C38002013402001A020800B0030AC;
    defparam PROG_MEM__D$n12.INIT_7 = 256'h0401100100180400601001820025010200845400C504615056A040012103100B;
    defparam PROG_MEM__D$n12.INIT_8 = 256'h420051021020020001002EA0219544EA041000000000D000000000000D0AD8BB;
    defparam PROG_MEM__D$n12.INIT_9 = 256'h0000000021820040051001C40020461000000000000001004000000400021000;
    defparam PROG_MEM__D$n12.INIT_A = 256'h0002102000100000000000000000000000040000000000001000040000000000;
    defparam PROG_MEM__D$n12.INIT_B = 256'h0204010000100000008000200000102000844841940AC084A8408C2840010030;
    defparam PROG_MEM__D$n12.INIT_C = 256'h0010821060000000205020832000022801010000000000001640050001421000;
    defparam PROG_MEM__D$n12.INIT_D = 256'h300010004002800B402818C3B0420430010018400010011000404000000C6080;
    defparam PROG_MEM__D$n12.INIT_E = 256'hC30A0232002B400C00D000003301B400818C38002013402001A020800B0030AC;
    defparam PROG_MEM__D$n12.INIT_F = 256'h0401100100180400601001820025010200845400C504615056A040012103100B;
    defparam PROG_MEM__D$n12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$n12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$n12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$n12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$n12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$n12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K USER_MEM__D$b12 (.WCLK(\CLK~O ), .RCLK(\CLK~O ), .WCLKE(n30807), 
            .WE(MEM_STORE), .RE(n50476), .WDATA({\SAVE_DATA[11] , \SAVE_DATA[10] , 
            \SAVE_DATA[9] , \SAVE_DATA[8] }), .WADDR({\SAVE_ADDRESS[9] , 
            \SAVE_ADDRESS[8] , \SAVE_ADDRESS[7] , \SAVE_ADDRESS[6] , \SAVE_ADDRESS[5] , 
            \SAVE_ADDRESS[4] , \SAVE_ADDRESS[3] , \SAVE_ADDRESS[2] , \SAVE_ADDRESS[1] , 
            \SAVE_ADDRESS[0] }), .RADDR({n1432, n1434, n1436, n1438, 
            n1440, n1442, n1444, n1446, n1448, n8}), .RDATA({\LOAD_DATA[11] , 
            \LOAD_DATA[10] , \LOAD_DATA[9] , \LOAD_DATA[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b0, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(234)
    defparam USER_MEM__D$b12.READ_WIDTH = 4;
    defparam USER_MEM__D$b12.WRITE_WIDTH = 4;
    defparam USER_MEM__D$b12.WCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$b12.WCLKE_POLARITY = 1'b1;
    defparam USER_MEM__D$b12.WE_POLARITY = 1'b1;
    defparam USER_MEM__D$b12.RCLK_POLARITY = 1'b1;
    defparam USER_MEM__D$b12.RE_POLARITY = 1'b0;
    defparam USER_MEM__D$b12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam USER_MEM__D$b12.OUTPUT_REG = 1'b0;
    defparam USER_MEM__D$b12.WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K PROG_MEM__D$m12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51742, 
            n51746})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h6106506902106106100103A88065133A800000000000DAAAAAAAAAAAA14111AD, INIT_1=256'h0102100610610214658230610618618000400000002000200000000000200630, INIT_2=256'h0000000002100000000000008000008000002000000000000000000211000200, INIT_3=256'h28420C010000400100400400000002800841840860C618618408408410000010, INIT_4=256'h8608608A81010660250000000200000720203001000A000108446505042908E0, INIT_5=256'h00220300B11710210290695B902106F402200010210200010800240200041161, INIT_6=256'h900B088314048200000003011000200014011000204250040140201033110052, INIT_7=256'hA03300A302028C0802302000001000060081060C2440840842002A0C0401082C, INIT_8=256'h6106506902106106100103A88065133A800000000000DAAAAAAAAAAAA14111AD, INIT_9=256'h0102100610610214658230610618618000400000002000200000000000200630, INIT_A=256'h0000000002100000000000008000008000002000000000000000000211000200, INIT_B=256'h28420C010000400100400400000002800841840860C618618408408410000010, INIT_C=256'h8608608A81010660250000000200000720203001000A000108446505042908E0, INIT_D=256'h00220300B11710210290695B902106F402200010210200010800240200041161, INIT_E=256'h900B088314048200000003011000200014011000204250040140201033110052, INIT_F=256'hA03300A302028C0802302000001000060081060C2440840842002A0C0401082C, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$m12.READ_WIDTH = 2;
    defparam PROG_MEM__D$m12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$m12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$m12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$m12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$m12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$m12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$m12.INIT_0 = 256'h6106506902106106100103A88065133A800000000000DAAAAAAAAAAAA14111AD;
    defparam PROG_MEM__D$m12.INIT_1 = 256'h0102100610610214658230610618618000400000002000200000000000200630;
    defparam PROG_MEM__D$m12.INIT_2 = 256'h0000000002100000000000008000008000002000000000000000000211000200;
    defparam PROG_MEM__D$m12.INIT_3 = 256'h28420C010000400100400400000002800841840860C618618408408410000010;
    defparam PROG_MEM__D$m12.INIT_4 = 256'h8608608A81010660250000000200000720203001000A000108446505042908E0;
    defparam PROG_MEM__D$m12.INIT_5 = 256'h00220300B11710210290695B902106F402200010210200010800240200041161;
    defparam PROG_MEM__D$m12.INIT_6 = 256'h900B088314048200000003011000200014011000204250040140201033110052;
    defparam PROG_MEM__D$m12.INIT_7 = 256'hA03300A302028C0802302000001000060081060C2440840842002A0C0401082C;
    defparam PROG_MEM__D$m12.INIT_8 = 256'h6106506902106106100103A88065133A800000000000DAAAAAAAAAAAA14111AD;
    defparam PROG_MEM__D$m12.INIT_9 = 256'h0102100610610214658230610618618000400000002000200000000000200630;
    defparam PROG_MEM__D$m12.INIT_A = 256'h0000000002100000000000008000008000002000000000000000000211000200;
    defparam PROG_MEM__D$m12.INIT_B = 256'h28420C010000400100400400000002800841840860C618618408408410000010;
    defparam PROG_MEM__D$m12.INIT_C = 256'h8608608A81010660250000000200000720203001000A000108446505042908E0;
    defparam PROG_MEM__D$m12.INIT_D = 256'h00220300B11710210290695B902106F402200010210200010800240200041161;
    defparam PROG_MEM__D$m12.INIT_E = 256'h900B088314048200000003011000200014011000204250040140201033110052;
    defparam PROG_MEM__D$m12.INIT_F = 256'hA03300A302028C0802302000001000060081060C2440840842002A0C0401082C;
    defparam PROG_MEM__D$m12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$m12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$m12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$m12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$m12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$m12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$l12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51750, 
            n51754})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0840840044840840800048EA0819048E200000000000EAAAAAAAAAAAA0104C64, INIT_1=256'h2000000084184084044084184004184010000000000000000000000000084084, INIT_2=256'h0840000000400000000000000040000400000000000000000000000000000000, INIT_3=256'h00451C000808008000002800000000000A38838818A782582182182180000000, INIT_4=256'h40AC10C028084104404010014000004010200000400200104090104000004294, INIT_5=256'h06004280000AC00300C0084E300A08F000000000000281010000000400018418, INIT_6=256'hE00C07417008C02C00000800AF00300808C4E300A0CC002002BC00C03486308E, INIT_7=256'h0000000C8200320800C82000500400020000505C09448005550008020002003F, INIT_8=256'h0840840044840840800048EA0819048E200000000000EAAAAAAAAAAAA0104C64, INIT_9=256'h2000000084184084044084184004184010000000000000000000000000084084, INIT_A=256'h0840000000400000000000000040000400000000000000000000000000000000, INIT_B=256'h00451C000808008000002800000000000A38838818A782582182182180000000, INIT_C=256'h40AC10C028084104404010014000004010200000400200104090104000004294, INIT_D=256'h06004280000AC00300C0084E300A08F000000000000281010000000400018418, INIT_E=256'hE00C07417008C02C00000800AF00300808C4E300A0CC002002BC00C03486308E, INIT_F=256'h0000000C8200320800C82000500400020000505C09448005550008020002003F, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$l12.READ_WIDTH = 2;
    defparam PROG_MEM__D$l12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$l12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$l12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$l12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$l12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$l12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$l12.INIT_0 = 256'h0840840044840840800048EA0819048E200000000000EAAAAAAAAAAAA0104C64;
    defparam PROG_MEM__D$l12.INIT_1 = 256'h2000000084184084044084184004184010000000000000000000000000084084;
    defparam PROG_MEM__D$l12.INIT_2 = 256'h0840000000400000000000000040000400000000000000000000000000000000;
    defparam PROG_MEM__D$l12.INIT_3 = 256'h00451C000808008000002800000000000A38838818A782582182182180000000;
    defparam PROG_MEM__D$l12.INIT_4 = 256'h40AC10C028084104404010014000004010200000400200104090104000004294;
    defparam PROG_MEM__D$l12.INIT_5 = 256'h06004280000AC00300C0084E300A08F000000000000281010000000400018418;
    defparam PROG_MEM__D$l12.INIT_6 = 256'hE00C07417008C02C00000800AF00300808C4E300A0CC002002BC00C03486308E;
    defparam PROG_MEM__D$l12.INIT_7 = 256'h0000000C8200320800C82000500400020000505C09448005550008020002003F;
    defparam PROG_MEM__D$l12.INIT_8 = 256'h0840840044840840800048EA0819048E200000000000EAAAAAAAAAAAA0104C64;
    defparam PROG_MEM__D$l12.INIT_9 = 256'h2000000084184084044084184004184010000000000000000000000000084084;
    defparam PROG_MEM__D$l12.INIT_A = 256'h0840000000400000000000000040000400000000000000000000000000000000;
    defparam PROG_MEM__D$l12.INIT_B = 256'h00451C000808008000002800000000000A38838818A782582182182180000000;
    defparam PROG_MEM__D$l12.INIT_C = 256'h40AC10C028084104404010014000004010200000400200104090104000004294;
    defparam PROG_MEM__D$l12.INIT_D = 256'h06004280000AC00300C0084E300A08F000000000000281010000000400018418;
    defparam PROG_MEM__D$l12.INIT_E = 256'hE00C07417008C02C00000800AF00300808C4E300A0CC002002BC00C03486308E;
    defparam PROG_MEM__D$l12.INIT_F = 256'h0000000C8200320800C82000500400020000505C09448005550008020002003F;
    defparam PROG_MEM__D$l12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$l12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$l12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$l12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$l12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$l12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$k12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51758, 
            n51762})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h840050A40840840848001238BA064123280000000000E0000000000001510544, INIT_1=256'h0008000060160851810020860840B60000000400020800000000000000800860, INIT_2=256'h0000000080000000800000001000002000021000000000041840004100040040, INIT_3=256'h2D0AD0002004036000400020801000C00D0200400818254A5201001020008008, INIT_4=256'h084083004086092080000A004208813C2D000820408C00110000850010210010, INIT_5=256'h10810080D40D508408408D8E40EC0FD002442C000000C0000040800040017004, INIT_6=256'h800820C001318300100000024100000C2486400480482018018800000084A14C, INIT_7=256'hA0800CA0D00A8340220D0080D900008900070840420270040210244900010012, INIT_8=256'h840050A40840840848001238BA064123280000000000E0000000000001510544, INIT_9=256'h0008000060160851810020860840B60000000400020800000000000000800860, INIT_A=256'h0000000080000000800000001000002000021000000000041840004100040040, INIT_B=256'h2D0AD0002004036000400020801000C00D0200400818254A5201001020008008, INIT_C=256'h084083004086092080000A004208813C2D000820408C00110000850010210010, INIT_D=256'h10810080D40D508408408D8E40EC0FD002442C000000C0000040800040017004, INIT_E=256'h800820C001318300100000024100000C2486400480482018018800000084A14C, INIT_F=256'hA0800CA0D00A8340220D0080D900008900070840420270040210244900010012, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$k12.READ_WIDTH = 2;
    defparam PROG_MEM__D$k12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$k12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$k12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$k12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$k12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$k12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$k12.INIT_0 = 256'h840050A40840840848001238BA064123280000000000E0000000000001510544;
    defparam PROG_MEM__D$k12.INIT_1 = 256'h0008000060160851810020860840B60000000400020800000000000000800860;
    defparam PROG_MEM__D$k12.INIT_2 = 256'h0000000080000000800000001000002000021000000000041840004100040040;
    defparam PROG_MEM__D$k12.INIT_3 = 256'h2D0AD0002004036000400020801000C00D0200400818254A5201001020008008;
    defparam PROG_MEM__D$k12.INIT_4 = 256'h084083004086092080000A004208813C2D000820408C00110000850010210010;
    defparam PROG_MEM__D$k12.INIT_5 = 256'h10810080D40D508408408D8E40EC0FD002442C000000C0000040800040017004;
    defparam PROG_MEM__D$k12.INIT_6 = 256'h800820C001318300100000024100000C2486400480482018018800000084A14C;
    defparam PROG_MEM__D$k12.INIT_7 = 256'hA0800CA0D00A8340220D0080D900008900070840420270040210244900010012;
    defparam PROG_MEM__D$k12.INIT_8 = 256'h840050A40840840848001238BA064123280000000000E0000000000001510544;
    defparam PROG_MEM__D$k12.INIT_9 = 256'h0008000060160851810020860840B60000000400020800000000000000800860;
    defparam PROG_MEM__D$k12.INIT_A = 256'h0000000080000000800000001000002000021000000000041840004100040040;
    defparam PROG_MEM__D$k12.INIT_B = 256'h2D0AD0002004036000400020801000C00D0200400818254A5201001020008008;
    defparam PROG_MEM__D$k12.INIT_C = 256'h084083004086092080000A004208813C2D000820408C00110000850010210010;
    defparam PROG_MEM__D$k12.INIT_D = 256'h10810080D40D508408408D8E40EC0FD002442C000000C0000040800040017004;
    defparam PROG_MEM__D$k12.INIT_E = 256'h800820C001318300100000024100000C2486400480482018018800000084A14C;
    defparam PROG_MEM__D$k12.INIT_F = 256'hA0800CA0D00A8340220D0080D900008900070840420270040210244900010012;
    defparam PROG_MEM__D$k12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$k12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$k12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$k12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$k12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$k12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$j12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51766, 
            n51770})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h01821860060821821800148CA4819148EA5C00000000C00000000000014F3AA8, INIT_1=256'h0000000618418614218200238218238008000010000010100000010000058218, INIT_2=256'h0000000000080000000002000000000000000000000000000800004002000000, INIT_3=256'h620038008000008000010400402000200960860960860CF89608608640000008, INIT_4=256'h4018118E00628228238008410000800804102810900000848298218208000608, INIT_5=256'h204028002089E80082FC19C8388D808800000000800000000000200200050860, INIT_6=256'h00021F116C100306120008009000002C49848108D008002003700000F5065104, INIT_7=256'h5000115040094100210400804004001000038108620208A0800880020802C034, INIT_8=256'h01821860060821821800148CA4819148EA5C00000000C00000000000014F3AA8, INIT_9=256'h0000000618418614218200238218238008000010000010100000010000058218, INIT_A=256'h0000000000080000000002000000000000000000000000000800004002000000, INIT_B=256'h620038008000008000010400402000200960860960860CF89608608640000008, INIT_C=256'h4018118E00628228238008410000800804102810900000848298218208000608, INIT_D=256'h204028002089E80082FC19C8388D808800000000800000000000200200050860, INIT_E=256'h00021F116C100306120008009000002C49848108D008002003700000F5065104, INIT_F=256'h5000115040094100210400804004001000038108620208A0800880020802C034, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$j12.READ_WIDTH = 2;
    defparam PROG_MEM__D$j12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$j12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$j12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$j12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$j12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$j12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$j12.INIT_0 = 256'h01821860060821821800148CA4819148EA5C00000000C00000000000014F3AA8;
    defparam PROG_MEM__D$j12.INIT_1 = 256'h0000000618418614218200238218238008000010000010100000010000058218;
    defparam PROG_MEM__D$j12.INIT_2 = 256'h0000000000080000000002000000000000000000000000000800004002000000;
    defparam PROG_MEM__D$j12.INIT_3 = 256'h620038008000008000010400402000200960860960860CF89608608640000008;
    defparam PROG_MEM__D$j12.INIT_4 = 256'h4018118E00628228238008410000800804102810900000848298218208000608;
    defparam PROG_MEM__D$j12.INIT_5 = 256'h204028002089E80082FC19C8388D808800000000800000000000200200050860;
    defparam PROG_MEM__D$j12.INIT_6 = 256'h00021F116C100306120008009000002C49848108D008002003700000F5065104;
    defparam PROG_MEM__D$j12.INIT_7 = 256'h5000115040094100210400804004001000038108620208A0800880020802C034;
    defparam PROG_MEM__D$j12.INIT_8 = 256'h01821860060821821800148CA4819148EA5C00000000C00000000000014F3AA8;
    defparam PROG_MEM__D$j12.INIT_9 = 256'h0000000618418614218200238218238008000010000010100000010000058218;
    defparam PROG_MEM__D$j12.INIT_A = 256'h0000000000080000000002000000000000000000000000000800004002000000;
    defparam PROG_MEM__D$j12.INIT_B = 256'h620038008000008000010400402000200960860960860CF89608608640000008;
    defparam PROG_MEM__D$j12.INIT_C = 256'h4018118E00628228238008410000800804102810900000848298218208000608;
    defparam PROG_MEM__D$j12.INIT_D = 256'h204028002089E80082FC19C8388D808800000000800000000000200200050860;
    defparam PROG_MEM__D$j12.INIT_E = 256'h00021F116C100306120008009000002C49848108D008002003700000F5065104;
    defparam PROG_MEM__D$j12.INIT_F = 256'h5000115040094100210400804004001000038108620208A0800880020802C034;
    defparam PROG_MEM__D$j12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$j12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$j12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$j12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$j12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$j12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$i12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51774, 
            n51778})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h9021021221121829020315231CA025123A4400000000EAAAAAAAAAAAA8D1A5CA, INIT_1=256'h0000000982D02180942142002106186000000008102130120001012000102102, INIT_2=256'h200032233001000000000000000000080D800000000002002002000010010000, INIT_3=256'h5001400200002080026010200000000804A840068848845842840840B0201003, INIT_4=256'h55C00041A85901001020060100011000224020224080808428001800A20C2D51, INIT_5=256'h500D00C0503D0310352B128D0193394000309012004004003100102000049002, INIT_6=256'h1C01042EC9000C21DE0C030310304200B050833830000000052040101AC0A121, INIT_7=256'h50422454100150400141001031015020800820069418001100809C2910028062, INIT_8=256'h9021021221121829020315231CA025123A4400000000EAAAAAAAAAAAA8D1A5CA, INIT_9=256'h0000000982D02180942142002106186000000008102130120001012000102102, INIT_A=256'h200032233001000000000000000000080D800000000002002002000010010000, INIT_B=256'h5001400200002080026010200000000804A840068848845842840840B0201003, INIT_C=256'h55C00041A85901001020060100011000224020224080808428001800A20C2D51, INIT_D=256'h500D00C0503D0310352B128D0193394000309012004004003100102000049002, INIT_E=256'h1C01042EC9000C21DE0C030310304200B050833830000000052040101AC0A121, INIT_F=256'h50422454100150400141001031015020800820069418001100809C2910028062, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$i12.READ_WIDTH = 2;
    defparam PROG_MEM__D$i12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$i12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$i12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$i12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$i12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$i12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$i12.INIT_0 = 256'h9021021221121829020315231CA025123A4400000000EAAAAAAAAAAAA8D1A5CA;
    defparam PROG_MEM__D$i12.INIT_1 = 256'h0000000982D02180942142002106186000000008102130120001012000102102;
    defparam PROG_MEM__D$i12.INIT_2 = 256'h200032233001000000000000000000080D800000000002002002000010010000;
    defparam PROG_MEM__D$i12.INIT_3 = 256'h5001400200002080026010200000000804A840068848845842840840B0201003;
    defparam PROG_MEM__D$i12.INIT_4 = 256'h55C00041A85901001020060100011000224020224080808428001800A20C2D51;
    defparam PROG_MEM__D$i12.INIT_5 = 256'h500D00C0503D0310352B128D0193394000309012004004003100102000049002;
    defparam PROG_MEM__D$i12.INIT_6 = 256'h1C01042EC9000C21DE0C030310304200B050833830000000052040101AC0A121;
    defparam PROG_MEM__D$i12.INIT_7 = 256'h50422454100150400141001031015020800820069418001100809C2910028062;
    defparam PROG_MEM__D$i12.INIT_8 = 256'h9021021221121829020315231CA025123A4400000000EAAAAAAAAAAAA8D1A5CA;
    defparam PROG_MEM__D$i12.INIT_9 = 256'h0000000982D02180942142002106186000000008102130120001012000102102;
    defparam PROG_MEM__D$i12.INIT_A = 256'h200032233001000000000000000000080D800000000002002002000010010000;
    defparam PROG_MEM__D$i12.INIT_B = 256'h5001400200002080026010200000000804A840068848845842840840B0201003;
    defparam PROG_MEM__D$i12.INIT_C = 256'h55C00041A85901001020060100011000224020224080808428001800A20C2D51;
    defparam PROG_MEM__D$i12.INIT_D = 256'h500D00C0503D0310352B128D0193394000309012004004003100102000049002;
    defparam PROG_MEM__D$i12.INIT_E = 256'h1C01042EC9000C21DE0C030310304200B050833830000000052040101AC0A121;
    defparam PROG_MEM__D$i12.INIT_F = 256'h50422454100150400141001031015020800820069418001100809C2910028062;
    defparam PROG_MEM__D$i12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$i12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$i12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$i12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$i12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$i12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$h12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51782, 
            n51786})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h86984D829861861860019448C1A889144E4404000000AAAAAAAAAAAAABC485C6, INIT_1=256'h02002008C18618A3840869A61865861000000000002B00000000000000861861, INIT_2=256'h0400000000010000000000000800000480800000000000000000000080000000, INIT_3=256'h860421000000104040400800000000200184180486D941941C41841840000041, INIT_4=256'h90208258848A08038200000000000245005000020C200006116A06A0888C9010, INIT_5=256'h000030002A1121C292713B7063025061000000200004000A0000080100002086, INIT_6=256'h3301BD04CC00081001000000100C00E4831301304200002000603030D40C4031, INIT_7=256'hA02208A0880A82202208808121A01021001001600400098082E8000008012044, INIT_8=256'h86984D829861861860019448C1A889144E4404000000AAAAAAAAAAAAABC485C6, INIT_9=256'h02002008C18618A3840869A61865861000000000002B00000000000000861861, INIT_A=256'h0400000000010000000000000800000480800000000000000000000080000000, INIT_B=256'h860421000000104040400800000000200184180486D941941C41841840000041, INIT_C=256'h90208258848A08038200000000000245005000020C200006116A06A0888C9010, INIT_D=256'h000030002A1121C292713B7063025061000000200004000A0000080100002086, INIT_E=256'h3301BD04CC00081001000000100C00E4831301304200002000603030D40C4031, INIT_F=256'hA02208A0880A82202208808121A01021001001600400098082E8000008012044, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$h12.READ_WIDTH = 2;
    defparam PROG_MEM__D$h12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$h12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$h12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$h12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$h12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$h12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$h12.INIT_0 = 256'h86984D829861861860019448C1A889144E4404000000AAAAAAAAAAAAABC485C6;
    defparam PROG_MEM__D$h12.INIT_1 = 256'h02002008C18618A3840869A61865861000000000002B00000000000000861861;
    defparam PROG_MEM__D$h12.INIT_2 = 256'h0400000000010000000000000800000480800000000000000000000080000000;
    defparam PROG_MEM__D$h12.INIT_3 = 256'h860421000000104040400800000000200184180486D941941C41841840000041;
    defparam PROG_MEM__D$h12.INIT_4 = 256'h90208258848A08038200000000000245005000020C200006116A06A0888C9010;
    defparam PROG_MEM__D$h12.INIT_5 = 256'h000030002A1121C292713B7063025061000000200004000A0000080100002086;
    defparam PROG_MEM__D$h12.INIT_6 = 256'h3301BD04CC00081001000000100C00E4831301304200002000603030D40C4031;
    defparam PROG_MEM__D$h12.INIT_7 = 256'hA02208A0880A82202208808121A01021001001600400098082E8000008012044;
    defparam PROG_MEM__D$h12.INIT_8 = 256'h86984D829861861860019448C1A889144E4404000000AAAAAAAAAAAAABC485C6;
    defparam PROG_MEM__D$h12.INIT_9 = 256'h02002008C18618A3840869A61865861000000000002B00000000000000861861;
    defparam PROG_MEM__D$h12.INIT_A = 256'h0400000000010000000000000800000480800000000000000000000080000000;
    defparam PROG_MEM__D$h12.INIT_B = 256'h860421000000104040400800000000200184180486D941941C41841840000041;
    defparam PROG_MEM__D$h12.INIT_C = 256'h90208258848A08038200000000000245005000020C200006116A06A0888C9010;
    defparam PROG_MEM__D$h12.INIT_D = 256'h000030002A1121C292713B7063025061000000200004000A0000080100002086;
    defparam PROG_MEM__D$h12.INIT_E = 256'h3301BD04CC00081001000000100C00E4831301304200002000603030D40C4031;
    defparam PROG_MEM__D$h12.INIT_F = 256'hA02208A0880A82202208808121A01021001001600400098082E8000008012044;
    defparam PROG_MEM__D$h12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$h12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$h12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$h12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$h12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$h12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$g12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51790, 
            n51794})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h50800845000840840A02645138EA225523080000000000000000000000515155, INIT_1=256'h0000000528408488418610108408408000000008000000400000000000408408, INIT_2=256'h0000800000040000000000000010001000000000000200000000000004001000, INIT_3=256'h4185080210000080A00000200000010C00210212210230A50A50210230000080, INIT_4=256'h000848044061064850A020024420008088400400008000108609008208318C1A, INIT_5=256'h4800A0C050F503C035A34A04C14A358300008820208000000400400000085860, INIT_6=256'h0580E24DCC020500020C00430038430C30A00E10E004300C7444400CE88CC024, INIT_7=256'h0840000A00C4280310A00C64C40000000001810141150010030949806A02C040, INIT_8=256'h50800845000840840A02645138EA225523080000000000000000000000515155, INIT_9=256'h0000000528408488418610108408408000000008000000400000000000408408, INIT_A=256'h0000800000040000000000000010001000000000000200000000000004001000, INIT_B=256'h4185080210000080A00000200000010C00210212210230A50A50210230000080, INIT_C=256'h000848044061064850A020024420008088400400008000108609008208318C1A, INIT_D=256'h4800A0C050F503C035A34A04C14A358300008820208000000400400000085860, INIT_E=256'h0580E24DCC020500020C00430038430C30A00E10E004300C7444400CE88CC024, INIT_F=256'h0840000A00C4280310A00C64C40000000001810141150010030949806A02C040, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$g12.READ_WIDTH = 2;
    defparam PROG_MEM__D$g12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$g12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$g12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$g12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$g12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$g12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$g12.INIT_0 = 256'h50800845000840840A02645138EA225523080000000000000000000000515155;
    defparam PROG_MEM__D$g12.INIT_1 = 256'h0000000528408488418610108408408000000008000000400000000000408408;
    defparam PROG_MEM__D$g12.INIT_2 = 256'h0000800000040000000000000010001000000000000200000000000004001000;
    defparam PROG_MEM__D$g12.INIT_3 = 256'h4185080210000080A00000200000010C00210212210230A50A50210230000080;
    defparam PROG_MEM__D$g12.INIT_4 = 256'h000848044061064850A020024420008088400400008000108609008208318C1A;
    defparam PROG_MEM__D$g12.INIT_5 = 256'h4800A0C050F503C035A34A04C14A358300008820208000000400400000085860;
    defparam PROG_MEM__D$g12.INIT_6 = 256'h0580E24DCC020500020C00430038430C30A00E10E004300C7444400CE88CC024;
    defparam PROG_MEM__D$g12.INIT_7 = 256'h0840000A00C4280310A00C64C40000000001810141150010030949806A02C040;
    defparam PROG_MEM__D$g12.INIT_8 = 256'h50800845000840840A02645138EA225523080000000000000000000000515155;
    defparam PROG_MEM__D$g12.INIT_9 = 256'h0000000528408488418610108408408000000008000000400000000000408408;
    defparam PROG_MEM__D$g12.INIT_A = 256'h0000800000040000000000000010001000000000000200000000000004001000;
    defparam PROG_MEM__D$g12.INIT_B = 256'h4185080210000080A00000200000010C00210212210230A50A50210230000080;
    defparam PROG_MEM__D$g12.INIT_C = 256'h000848044061064850A020024420008088400400008000108609008208318C1A;
    defparam PROG_MEM__D$g12.INIT_D = 256'h4800A0C050F503C035A34A04C14A358300008820208000000400400000085860;
    defparam PROG_MEM__D$g12.INIT_E = 256'h0580E24DCC020500020C00430038430C30A00E10E004300C7444400CE88CC024;
    defparam PROG_MEM__D$g12.INIT_F = 256'h0840000A00C4280310A00C64C40000000001810141150010030949806A02C040;
    defparam PROG_MEM__D$g12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$g12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$g12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$g12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$g12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$g12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$f12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51798, 
            n51802})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0841841B4004184124009854BF3A899548800000000020000000000003024F98, INIT_1=256'h00008401241841861860800B4186183000000000010000812000001040184084, INIT_2=256'h08008840000000000000000000000000000020000000002000000040840A0080, INIT_3=256'h11010600000420B000006B00800000000610610410610754E106106100000000, INIT_4=256'h618318000F2143041050000804A209C0804800008820C04801A51242A56850B0, INIT_5=256'hC04000004A40A4884CBD3D408D0A40840208040201401090C080000008008628, INIT_6=256'h0620F4E05400EC1909040800000C00D081480080400800300040E00344090408, INIT_7=256'h002C0800300000C00003000808008910800805A206A041721A31035005030C84, INIT_8=256'h0841841B4004184124009854BF3A899548800000000020000000000003024F98, INIT_9=256'h00008401241841861860800B4186183000000000010000812000001040184084, INIT_A=256'h08008840000000000000000000000000000020000000002000000040840A0080, INIT_B=256'h11010600000420B000006B00800000000610610410610754E106106100000000, INIT_C=256'h618318000F2143041050000804A209C0804800008820C04801A51242A56850B0, INIT_D=256'hC04000004A40A4884CBD3D408D0A40840208040201401090C080000008008628, INIT_E=256'h0620F4E05400EC1909040800000C00D081480080400800300040E00344090408, INIT_F=256'h002C0800300000C00003000808008910800805A206A041721A31035005030C84, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$f12.READ_WIDTH = 2;
    defparam PROG_MEM__D$f12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$f12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$f12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$f12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$f12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$f12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$f12.INIT_0 = 256'h0841841B4004184124009854BF3A899548800000000020000000000003024F98;
    defparam PROG_MEM__D$f12.INIT_1 = 256'h00008401241841861860800B4186183000000000010000812000001040184084;
    defparam PROG_MEM__D$f12.INIT_2 = 256'h08008840000000000000000000000000000020000000002000000040840A0080;
    defparam PROG_MEM__D$f12.INIT_3 = 256'h11010600000420B000006B00800000000610610410610754E106106100000000;
    defparam PROG_MEM__D$f12.INIT_4 = 256'h618318000F2143041050000804A209C0804800008820C04801A51242A56850B0;
    defparam PROG_MEM__D$f12.INIT_5 = 256'hC04000004A40A4884CBD3D408D0A40840208040201401090C080000008008628;
    defparam PROG_MEM__D$f12.INIT_6 = 256'h0620F4E05400EC1909040800000C00D081480080400800300040E00344090408;
    defparam PROG_MEM__D$f12.INIT_7 = 256'h002C0800300000C00003000808008910800805A206A041721A31035005030C84;
    defparam PROG_MEM__D$f12.INIT_8 = 256'h0841841B4004184124009854BF3A899548800000000020000000000003024F98;
    defparam PROG_MEM__D$f12.INIT_9 = 256'h00008401241841861860800B4186183000000000010000812000001040184084;
    defparam PROG_MEM__D$f12.INIT_A = 256'h08008840000000000000000000000000000020000000002000000040840A0080;
    defparam PROG_MEM__D$f12.INIT_B = 256'h11010600000420B000006B00800000000610610410610754E106106100000000;
    defparam PROG_MEM__D$f12.INIT_C = 256'h618318000F2143041050000804A209C0804800008820C04801A51242A56850B0;
    defparam PROG_MEM__D$f12.INIT_D = 256'hC04000004A40A4884CBD3D408D0A40840208040201401090C080000008008628;
    defparam PROG_MEM__D$f12.INIT_E = 256'h0620F4E05400EC1909040800000C00D081480080400800300040E00344090408;
    defparam PROG_MEM__D$f12.INIT_F = 256'h002C0800300000C00003000808008910800805A206A041721A31035005030C84;
    defparam PROG_MEM__D$f12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$f12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$f12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$f12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$f12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$f12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$e12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51806, 
            n51810})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h821021001921021020020655008EA0255200000000004AAAAAAAAAAAAA1A59DD, INIT_1=256'h0000100821821021C01061821021061000004018000001010000000000041421, INIT_2=256'h20000000101000000000C0000044000010000000000000000000000000000400, INIT_3=256'h0A0060000000104000000900000000000086282086A8609E8860860CE0000001, INIT_4=256'h30610009600E10900400100800A10818000000002C0080129010C21440120504, INIT_5=256'h60C6000000C6300020B14814014B041000000000008087001801000100024182, INIT_6=256'h43003BC480730400728401002100002B138118108003000032848000B4E10610, INIT_7=256'h0008010100300400C010030180000910004408551220214698E91C19200300BC, INIT_8=256'h821021001921021020020655008EA0255200000000004AAAAAAAAAAAAA1A59DD, INIT_9=256'h0000100821821021C01061821021061000004018000001010000000000041421, INIT_A=256'h20000000101000000000C0000044000010000000000000000000000000000400, INIT_B=256'h0A0060000000104000000900000000000086282086A8609E8860860CE0000001, INIT_C=256'h30610009600E10900400100800A10818000000002C0080129010C21440120504, INIT_D=256'h60C6000000C6300020B14814014B041000000000008087001801000100024182, INIT_E=256'h43003BC480730400728401002100002B138118108003000032848000B4E10610, INIT_F=256'h0008010100300400C010030180000910004408551220214698E91C19200300BC, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$e12.READ_WIDTH = 2;
    defparam PROG_MEM__D$e12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$e12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$e12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$e12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$e12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$e12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$e12.INIT_0 = 256'h821021001921021020020655008EA0255200000000004AAAAAAAAAAAAA1A59DD;
    defparam PROG_MEM__D$e12.INIT_1 = 256'h0000100821821021C01061821021061000004018000001010000000000041421;
    defparam PROG_MEM__D$e12.INIT_2 = 256'h20000000101000000000C0000044000010000000000000000000000000000400;
    defparam PROG_MEM__D$e12.INIT_3 = 256'h0A0060000000104000000900000000000086282086A8609E8860860CE0000001;
    defparam PROG_MEM__D$e12.INIT_4 = 256'h30610009600E10900400100800A10818000000002C0080129010C21440120504;
    defparam PROG_MEM__D$e12.INIT_5 = 256'h60C6000000C6300020B14814014B041000000000008087001801000100024182;
    defparam PROG_MEM__D$e12.INIT_6 = 256'h43003BC480730400728401002100002B138118108003000032848000B4E10610;
    defparam PROG_MEM__D$e12.INIT_7 = 256'h0008010100300400C010030180000910004408551220214698E91C19200300BC;
    defparam PROG_MEM__D$e12.INIT_8 = 256'h821021001921021020020655008EA0255200000000004AAAAAAAAAAAAA1A59DD;
    defparam PROG_MEM__D$e12.INIT_9 = 256'h0000100821821021C01061821021061000004018000001010000000000041421;
    defparam PROG_MEM__D$e12.INIT_A = 256'h20000000101000000000C0000044000010000000000000000000000000000400;
    defparam PROG_MEM__D$e12.INIT_B = 256'h0A0060000000104000000900000000000086282086A8609E8860860CE0000001;
    defparam PROG_MEM__D$e12.INIT_C = 256'h30610009600E10900400100800A10818000000002C0080129010C21440120504;
    defparam PROG_MEM__D$e12.INIT_D = 256'h60C6000000C6300020B14814014B041000000000008087001801000100024182;
    defparam PROG_MEM__D$e12.INIT_E = 256'h43003BC480730400728401002100002B138118108003000032848000B4E10610;
    defparam PROG_MEM__D$e12.INIT_F = 256'h0008010100300400C010030180000910004408551220214698E91C19200300BC;
    defparam PROG_MEM__D$e12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$e12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$e12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$e12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$e12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$e12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$d12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51814, 
            n51818})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'hE1060069861061060002819541238899548C00000000EAAAAAAAAAAAAA88EA82, INIT_1=256'h0000100E08610690C30684E40610658000800000000403900000000400650614, INIT_2=256'h0020020210020000010000000400000000408400004000040020000800240240, INIT_3=256'h6046C4000800200000C00248000000800C4084A84084084C9408408400202000, INIT_4=256'h061C20C450440A122A2010000260000648040A00200400210204E90444410296, INIT_5=256'h012820002106102107123107D06D025000200400230030008020000200023800, INIT_6=256'hA080040A2674870AA04804204000005831025824010800000340000050812070, INIT_7=256'h0101020000200000800002212010500040099880115680094010268110010834, INIT_8=256'hE1060069861061060002819541238899548C00000000EAAAAAAAAAAAAA88EA82, INIT_9=256'h0000100E08610690C30684E40610658000800000000403900000000400650614, INIT_A=256'h0020020210020000010000000400000000408400004000040020000800240240, INIT_B=256'h6046C4000800200000C00248000000800C4084A84084084C9408408400202000, INIT_C=256'h061C20C450440A122A2010000260000648040A00200400210204E90444410296, INIT_D=256'h012820002106102107123107D06D025000200400230030008020000200023800, INIT_E=256'hA080040A2674870AA04804204000005831025824010800000340000050812070, INIT_F=256'h0101020000200000800002212010500040099880115680094010268110010834, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$d12.READ_WIDTH = 2;
    defparam PROG_MEM__D$d12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$d12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$d12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$d12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$d12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$d12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$d12.INIT_0 = 256'hE1060069861061060002819541238899548C00000000EAAAAAAAAAAAAA88EA82;
    defparam PROG_MEM__D$d12.INIT_1 = 256'h0000100E08610690C30684E40610658000800000000403900000000400650614;
    defparam PROG_MEM__D$d12.INIT_2 = 256'h0020020210020000010000000400000000408400004000040020000800240240;
    defparam PROG_MEM__D$d12.INIT_3 = 256'h6046C4000800200000C00248000000800C4084A84084084C9408408400202000;
    defparam PROG_MEM__D$d12.INIT_4 = 256'h061C20C450440A122A2010000260000648040A00200400210204E90444410296;
    defparam PROG_MEM__D$d12.INIT_5 = 256'h012820002106102107123107D06D025000200400230030008020000200023800;
    defparam PROG_MEM__D$d12.INIT_6 = 256'hA080040A2674870AA04804204000005831025824010800000340000050812070;
    defparam PROG_MEM__D$d12.INIT_7 = 256'h0101020000200000800002212010500040099880115680094010268110010834;
    defparam PROG_MEM__D$d12.INIT_8 = 256'hE1060069861061060002819541238899548C00000000EAAAAAAAAAAAAA88EA82;
    defparam PROG_MEM__D$d12.INIT_9 = 256'h0000100E08610690C30684E40610658000800000000403900000000400650614;
    defparam PROG_MEM__D$d12.INIT_A = 256'h0020020210020000010000000400000000408400004000040020000800240240;
    defparam PROG_MEM__D$d12.INIT_B = 256'h6046C4000800200000C00248000000800C4084A84084084C9408408400202000;
    defparam PROG_MEM__D$d12.INIT_C = 256'h061C20C450440A122A2010000260000648040A00200400210204E90444410296;
    defparam PROG_MEM__D$d12.INIT_D = 256'h012820002106102107123107D06D025000200400230030008020000200023800;
    defparam PROG_MEM__D$d12.INIT_E = 256'hA080040A2674870AA04804204000005831025824010800000340000050812070;
    defparam PROG_MEM__D$d12.INIT_F = 256'h0101020000200000800002212010500040099880115680094010268110010834;
    defparam PROG_MEM__D$d12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$d12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$d12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$d12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$d12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$d12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$c12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51822, 
            n51826})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0860860860820860860222655148C20655140000000040000000000000544115, INIT_1=256'h0000100086181086182006186086082000004000000004000000000000086086, INIT_2=256'h0000000020C00000000000000010000000000000000000000000000000200000, INIT_3=256'h002004000008304010800000100000080A380142182182382382182190000042, INIT_4=256'h208485A1043001000260000008000840440A0144200240086582080284004080, INIT_5=256'h00E40000002236002A36003AC28FF0D30200009000000080048220A000018A98, INIT_6=256'h4000B8C0005F0230C38C0400634000E30001AC58C10F1020028404028D0424B1, INIT_7=256'h005002005080014200050810400010200010430208600290210208A10000403C, INIT_8=256'h0860860860820860860222655148C20655140000000040000000000000544115, INIT_9=256'h0000100086181086182006186086082000004000000004000000000000086086, INIT_A=256'h0000000020C00000000000000010000000000000000000000000000000200000, INIT_B=256'h002004000008304010800000100000080A380142182182382382182190000042, INIT_C=256'h208485A1043001000260000008000840440A0144200240086582080284004080, INIT_D=256'h00E40000002236002A36003AC28FF0D30200009000000080048220A000018A98, INIT_E=256'h4000B8C0005F0230C38C0400634000E30001AC58C10F1020028404028D0424B1, INIT_F=256'h005002005080014200050810400010200010430208600290210208A10000403C, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$c12.READ_WIDTH = 2;
    defparam PROG_MEM__D$c12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$c12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$c12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$c12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$c12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$c12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$c12.INIT_0 = 256'h0860860860820860860222655148C20655140000000040000000000000544115;
    defparam PROG_MEM__D$c12.INIT_1 = 256'h0000100086181086182006186086082000004000000004000000000000086086;
    defparam PROG_MEM__D$c12.INIT_2 = 256'h0000000020C00000000000000010000000000000000000000000000000200000;
    defparam PROG_MEM__D$c12.INIT_3 = 256'h002004000008304010800000100000080A380142182182382382182190000042;
    defparam PROG_MEM__D$c12.INIT_4 = 256'h208485A1043001000260000008000840440A0144200240086582080284004080;
    defparam PROG_MEM__D$c12.INIT_5 = 256'h00E40000002236002A36003AC28FF0D30200009000000080048220A000018A98;
    defparam PROG_MEM__D$c12.INIT_6 = 256'h4000B8C0005F0230C38C0400634000E30001AC58C10F1020028404028D0424B1;
    defparam PROG_MEM__D$c12.INIT_7 = 256'h005002005080014200050810400010200010430208600290210208A10000403C;
    defparam PROG_MEM__D$c12.INIT_8 = 256'h0860860860820860860222655148C20655140000000040000000000000544115;
    defparam PROG_MEM__D$c12.INIT_9 = 256'h0000100086181086182006186086082000004000000004000000000000086086;
    defparam PROG_MEM__D$c12.INIT_A = 256'h0000000020C00000000000000010000000000000000000000000000000200000;
    defparam PROG_MEM__D$c12.INIT_B = 256'h002004000008304010800000100000080A380142182182382382182190000042;
    defparam PROG_MEM__D$c12.INIT_C = 256'h208485A1043001000260000008000840440A0144200240086582080284004080;
    defparam PROG_MEM__D$c12.INIT_D = 256'h00E40000002236002A36003AC28FF0D30200009000000080048220A000018A98;
    defparam PROG_MEM__D$c12.INIT_E = 256'h4000B8C0005F0230C38C0400634000E30001AC58C10F1020028404028D0424B1;
    defparam PROG_MEM__D$c12.INIT_F = 256'h005002005080014200050810400010200010430208600290210208A10000403C;
    defparam PROG_MEM__D$c12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$c12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$c12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$c12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$c12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$c12.WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K PROG_MEM__D$12 (.WCLK(1'b0), .RCLK(\CLK~O ), .WCLKE(1'b0), 
            .WE(1'b0), .RE(1'b1), .WADDR({11'b00000000000}), .RADDR({\PC[10] , 
            \PC[9] , \PC[8] , \PC[7] , \PC[6] , \PC[5] , \PC[4] , 
            \PC[3] , \PC[2] , \PC[1] , \PC[0]__I }), .RDATA({n51838, 
            n51842})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h21821A21811021800800420641148C206500000000001AAAAAAAAAAAA892A288, INIT_1=256'h000008063802A218238619218618238000000000012040000100000000218018, INIT_2=256'h0000000000000000000000000000002000100000002000000000000000000000, INIT_3=256'h21213B000000000030302408000008300861861861C618719618619630000008, INIT_4=256'h020A428201208630418004000200880A1001000221000001821000B223008142, INIT_5=256'hC014008000881E31A81D01814A82E3C90000001000A008048000091800040842, INIT_6=256'h554430400A909B304004080080411081000018080030202C02050C460DC04800, INIT_7=256'h51240050298140A6050298158400014080612D1260A00308248400A01102C030, INIT_8=256'h21821A21811021800800420641148C206500000000001AAAAAAAAAAAA892A288, INIT_9=256'h000008063802A218238619218618238000000000012040000100000000218018, INIT_A=256'h0000000000000000000000000000002000100000002000000000000000000000, INIT_B=256'h21213B000000000030302408000008300861861861C618719618619630000008, INIT_C=256'h020A428201208630418004000200880A1001000221000001821000B223008142, INIT_D=256'hC014008000881E31A81D01814A82E3C90000001000A008048000091800040842, INIT_E=256'h554430400A909B304004080080411081000018080030202C02050C460DC04800, INIT_F=256'h51240050298140A6050298158400014080612D1260A00308248400A01102C030, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(47)
    defparam PROG_MEM__D$12.READ_WIDTH = 2;
    defparam PROG_MEM__D$12.WRITE_WIDTH = 2;
    defparam PROG_MEM__D$12.WCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$12.WCLKE_POLARITY = 1'b1;
    defparam PROG_MEM__D$12.WE_POLARITY = 1'b1;
    defparam PROG_MEM__D$12.RCLK_POLARITY = 1'b1;
    defparam PROG_MEM__D$12.RE_POLARITY = 1'b1;
    defparam PROG_MEM__D$12.INIT_0 = 256'h21821A21811021800800420641148C206500000000001AAAAAAAAAAAA892A288;
    defparam PROG_MEM__D$12.INIT_1 = 256'h000008063802A218238619218618238000000000012040000100000000218018;
    defparam PROG_MEM__D$12.INIT_2 = 256'h0000000000000000000000000000002000100000002000000000000000000000;
    defparam PROG_MEM__D$12.INIT_3 = 256'h21213B000000000030302408000008300861861861C618719618619630000008;
    defparam PROG_MEM__D$12.INIT_4 = 256'h020A428201208630418004000200880A1001000221000001821000B223008142;
    defparam PROG_MEM__D$12.INIT_5 = 256'hC014008000881E31A81D01814A82E3C90000001000A008048000091800040842;
    defparam PROG_MEM__D$12.INIT_6 = 256'h554430400A909B304004080080411081000018080030202C02050C460DC04800;
    defparam PROG_MEM__D$12.INIT_7 = 256'h51240050298140A6050298158400014080612D1260A00308248400A01102C030;
    defparam PROG_MEM__D$12.INIT_8 = 256'h21821A21811021800800420641148C206500000000001AAAAAAAAAAAA892A288;
    defparam PROG_MEM__D$12.INIT_9 = 256'h000008063802A218238619218618238000000000012040000100000000218018;
    defparam PROG_MEM__D$12.INIT_A = 256'h0000000000000000000000000000002000100000002000000000000000000000;
    defparam PROG_MEM__D$12.INIT_B = 256'h21213B000000000030302408000008300861861861C618719618619630000008;
    defparam PROG_MEM__D$12.INIT_C = 256'h020A428201208630418004000200880A1001000221000001821000B223008142;
    defparam PROG_MEM__D$12.INIT_D = 256'hC014008000881E31A81D01814A82E3C90000001000A008048000091800040842;
    defparam PROG_MEM__D$12.INIT_E = 256'h554430400A909B304004080080411081000018080030202C02050C460DC04800;
    defparam PROG_MEM__D$12.INIT_F = 256'h51240050298140A6050298158400014080612D1260A00308248400A01102C030;
    defparam PROG_MEM__D$12.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$12.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$12.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$12.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam PROG_MEM__D$12.OUTPUT_REG = 1'b0;
    defparam PROG_MEM__D$12.WRITE_MODE = "READ_UNKNOWN";
    EFX_LUT4 LUT__4495 (.I0(\XI[1][26] ), .I1(\XI[0][26] ), .I2(n2953), 
            .I3(n2954), .O(n2955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4495.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4496 (.I0(\XI[3][26] ), .I1(\XI[2][26] ), .I2(n2954), 
            .I3(n2953), .O(n2956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4496.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4497 (.I0(\XI[7][26] ), .I1(\XI[5][26] ), .I2(n2954), 
            .I3(n2953), .O(n2957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4497.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4498 (.I0(\XI[6][26] ), .I1(\XI[4][26] ), .I2(n2954), 
            .I3(n2957), .O(n2958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4498.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4499 (.I0(STAGE2_EN), .I1(n51762), .O(n2959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4499.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4500 (.I0(n2956), .I1(n2955), .I2(n2958), .I3(n2959), 
            .O(n2960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__4500.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__4501 (.I0(\XI[9][26] ), .I1(\XI[8][26] ), .I2(n2953), 
            .I3(n2954), .O(n2961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4501.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4502 (.I0(\XI[11][26] ), .I1(\XI[10][26] ), .I2(n2954), 
            .I3(n2953), .O(n2962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4502.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4503 (.I0(\XI[15][26] ), .I1(\XI[13][26] ), .I2(n2954), 
            .I3(n2953), .O(n2963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4503.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4504 (.I0(\XI[14][26] ), .I1(\XI[12][26] ), .I2(n2954), 
            .I3(n2963), .O(n2964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4504.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4505 (.I0(n2962), .I1(n2961), .I2(n2964), .I3(n2959), 
            .O(n2965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__4505.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__4506 (.I0(STAGE2_EN), .I1(n51754), .O(n2966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4506.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4507 (.I0(STAGE2_EN), .I1(n51758), .O(n2967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4507.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4508 (.I0(n2965), .I1(n2960), .I2(n2966), .I3(n2967), 
            .O(n2968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4508.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4509 (.I0(\XI[29][26] ), .I1(\XI[28][26] ), .I2(n2953), 
            .I3(n2954), .O(n2969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4509.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4510 (.I0(\XI[31][26] ), .I1(\XI[30][26] ), .I2(n2954), 
            .I3(n2953), .O(n2970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4510.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4511 (.I0(\XI[27][26] ), .I1(\XI[25][26] ), .I2(n2954), 
            .I3(n2953), .O(n2971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4511.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4512 (.I0(\XI[26][26] ), .I1(\XI[24][26] ), .I2(n2954), 
            .I3(n2971), .O(n2972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4512.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4513 (.I0(n2970), .I1(n2969), .I2(n2972), .I3(n2959), 
            .O(n2973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4513.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4514 (.I0(\XI[23][26] ), .I1(\XI[22][26] ), .I2(n2954), 
            .I3(n2953), .O(n2974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4514.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4515 (.I0(\XI[21][26] ), .I1(\XI[20][26] ), .I2(n2953), 
            .I3(n2954), .O(n2975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4515.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4516 (.I0(\XI[19][26] ), .I1(\XI[17][26] ), .I2(n2954), 
            .I3(n2953), .O(n2976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4516.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4517 (.I0(\XI[18][26] ), .I1(\XI[16][26] ), .I2(n2954), 
            .I3(n2976), .O(n2977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4517.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4518 (.I0(n2975), .I1(n2974), .I2(n2977), .I3(n2959), 
            .O(n2978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4518.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4519 (.I0(n2978), .I1(n2973), .I2(n2967), .I3(n2966), 
            .O(n2979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__4519.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__4520 (.I0(n51834), .I1(n51826), .I2(STAGE2_EN), .I3(n51830), 
            .O(n2980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__4520.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__4521 (.I0(n2980), .I1(n51842), .O(n2981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4521.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4522 (.I0(n51834), .I1(STAGE2_EN), .O(n2982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4522.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4523 (.I0(n51838), .I1(n51842), .I2(n2982), .O(n2983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4523.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4524 (.I0(n51834), .I1(n51842), .I2(n51838), .I3(STAGE2_EN), 
            .O(n2984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__4524.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__4525 (.I0(n2983), .I1(n2980), .I2(n2984), .O(n2985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__4525.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__4526 (.I0(STAGE2_EN), .I1(n51826), .O(n2986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4526.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4527 (.I0(n2985), .I1(n2981), .I2(n2986), .O(n2987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__4527.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__4528 (.I0(\PC[26] ), .I1(n51726), .I2(n51838), .O(n2988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4528.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4529 (.I0(n51842), .I1(n51838), .O(n2989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__4529.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__4530 (.I0(n2989), .I1(n51726), .I2(n51830), .I3(STAGE2_EN), 
            .O(n2990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__4530.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__4531 (.I0(n2984), .I1(n2990), .O(n2991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4531.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4532 (.I0(n2983), .I1(\PC[26] ), .I2(n2991), .O(n2992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__4532.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__4533 (.I0(n2981), .I1(n2988), .I2(n2992), .I3(n2986), 
            .O(n2993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__4533.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__4534 (.I0(n2979), .I1(n2968), .I2(n2987), .I3(n2993), 
            .O(n500_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff */ ;
    defparam LUT__4534.LUTMASK = 16'h10ff;
    EFX_LUT4 LUT__4535 (.I0(STAGE2_EN), .I1(n221), .O(n30664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4535.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4536 (.I0(\XII[16][4] ), .I1(\XII[18][4] ), .I2(n51766), 
            .O(n2994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4536.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4537 (.I0(\XII[17][4] ), .I1(\XII[19][4] ), .I2(n51766), 
            .O(n2995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4537.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4538 (.I0(n2995), .I1(n2994), .I2(n2959), .I3(n2954), 
            .O(n2996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4538.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4539 (.I0(\XII[20][4] ), .I1(\XII[22][4] ), .I2(n51766), 
            .O(n2997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4539.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4540 (.I0(\XII[21][4] ), .I1(\XII[23][4] ), .I2(n51766), 
            .O(n2998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4540.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4541 (.I0(n2998), .I1(n2997), .I2(n2954), .I3(n2959), 
            .O(n2999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4541.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4542 (.I0(n2996), .I1(n2999), .I2(n2967), .O(n3000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__4542.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__4543 (.I0(\XII[28][4] ), .I1(\XII[30][4] ), .I2(n51766), 
            .O(n3001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4543.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4544 (.I0(\XII[29][4] ), .I1(\XII[31][4] ), .I2(n51766), 
            .O(n3002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4544.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4545 (.I0(n3002), .I1(n3001), .I2(n2954), .I3(n2959), 
            .O(n3003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4545.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4546 (.I0(\XII[24][4] ), .I1(\XII[26][4] ), .I2(n51766), 
            .O(n3004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4546.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4547 (.I0(\XII[25][4] ), .I1(\XII[27][4] ), .I2(n51766), 
            .O(n3005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4547.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4548 (.I0(n3005), .I1(n3004), .I2(n2959), .I3(n2954), 
            .O(n3006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4548.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4549 (.I0(n3006), .I1(n3003), .I2(n2967), .I3(n2966), 
            .O(n3007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__4549.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__4556 (.I0(n3013), .I1(n3010), .I2(n2959), .I3(n2967), 
            .O(n3014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4556.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4557 (.I0(\XII[0][4] ), .I1(\XII[2][4] ), .I2(n51766), 
            .O(n3015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__4557.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__4558 (.I0(\XII[1][4] ), .I1(\XII[3][4] ), .I2(n51766), 
            .O(n3016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__4558.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__4559 (.I0(n3016), .I1(n3015), .I2(n2959), .I3(n2954), 
            .O(n3017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4559.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4560 (.I0(\XII[4][4] ), .I1(\XII[6][4] ), .I2(n51766), 
            .O(n3018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__4560.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__4561 (.I0(\XII[5][4] ), .I1(\XII[7][4] ), .I2(n51766), 
            .O(n3019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__4561.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__4562 (.I0(n3019), .I1(n3018), .I2(n2954), .I3(n2959), 
            .O(n3020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4562.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4563 (.I0(n3020), .I1(n2967), .I2(n3017), .I3(n2966), 
            .O(n3021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__4563.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__4564 (.I0(n3014), .I1(n3021), .I2(n3000), .I3(n3007), 
            .O(n3022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__4564.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__4565 (.I0(n2983), .I1(n3022), .I2(n51830), .I3(n2984), 
            .O(n3023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heee0 */ ;
    defparam LUT__4565.LUTMASK = 16'heee0;
    EFX_LUT4 LUT__4566 (.I0(\PC[4] ), .I1(n51834), .I2(n51754), .I3(n51842), 
            .O(n3024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__4566.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__4567 (.I0(n51830), .I1(n51838), .I2(n3024), .I3(n51826), 
            .O(n3025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__4567.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__4568 (.I0(n51834), .I1(n51830), .I2(STAGE2_EN), .I3(n51838), 
            .O(n3026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__4568.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__4569 (.I0(\PC[4] ), .I1(n51754), .I2(n3026), .O(n3027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4569.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4570 (.I0(n51834), .I1(n51830), .I2(STAGE2_EN), .O(n3028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4570.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4571 (.I0(n3028), .I1(n51842), .O(n3029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4571.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4572 (.I0(n3022), .I1(n3027), .I2(n3029), .I3(n2986), 
            .O(n3030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__4572.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__4573 (.I0(n3023), .I1(n3025), .I2(STAGE2_EN), .I3(n3030), 
            .O(n522_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__4573.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__4574 (.I0(\XII[5][3] ), .I1(\XII[4][3] ), .I2(n2953), 
            .I3(n2954), .O(n3031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4574.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4575 (.I0(\XII[7][3] ), .I1(\XII[6][3] ), .I2(n2954), 
            .I3(n2953), .O(n3032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4575.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4576 (.I0(\XII[1][3] ), .I1(\XII[0][3] ), .I2(STAGE2_EN), 
            .I3(n51770), .O(n3033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333 */ ;
    defparam LUT__4576.LUTMASK = 16'h5333;
    EFX_LUT4 LUT__4577 (.I0(\XII[2][3] ), .I1(\XII[3][3] ), .I2(n51770), 
            .O(n3034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4577.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4578 (.I0(n3034), .I1(n3033), .I2(n2953), .O(n3035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__4578.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__4579 (.I0(n3032), .I1(n3031), .I2(n3035), .I3(n2959), 
            .O(n3036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4579.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4580 (.I0(\XII[13][3] ), .I1(\XII[12][3] ), .I2(n2953), 
            .I3(n2954), .O(n3037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4580.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4581 (.I0(\XII[15][3] ), .I1(\XII[14][3] ), .I2(n2954), 
            .I3(n2953), .O(n3038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4581.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4585 (.I0(n3038), .I1(n3037), .I2(n3041), .I3(n2959), 
            .O(n3042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4585.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4586 (.I0(n3042), .I1(n3036), .I2(n2966), .I3(n2967), 
            .O(n3043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4586.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4587 (.I0(\XII[26][3] ), .I1(\XII[27][3] ), .I2(n51770), 
            .O(n3044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4587.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4588 (.I0(\XII[24][3] ), .I1(\XII[25][3] ), .I2(n51770), 
            .O(n3045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4588.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4589 (.I0(n3044), .I1(n3045), .I2(n2967), .I3(n2953), 
            .O(n3046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4589.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4590 (.I0(\XII[21][3] ), .I1(\XII[20][3] ), .I2(n2953), 
            .I3(n2954), .O(n3047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4590.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4591 (.I0(\XII[23][3] ), .I1(\XII[22][3] ), .I2(n51770), 
            .O(n3048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4591.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4592 (.I0(n3048), .I1(n3046), .I2(n3047), .I3(n2967), 
            .O(n3049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h330e */ ;
    defparam LUT__4592.LUTMASK = 16'h330e;
    EFX_LUT4 LUT__4593 (.I0(\XII[28][3] ), .I1(\XII[29][3] ), .I2(n51770), 
            .O(n3050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4593.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4594 (.I0(\XII[30][3] ), .I1(\XII[31][3] ), .I2(n51770), 
            .O(n3051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4594.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4595 (.I0(n3051), .I1(n3050), .I2(n2953), .I3(n2959), 
            .O(n3052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4595.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4596 (.I0(\XII[16][3] ), .I1(\XII[17][3] ), .I2(n51770), 
            .O(n3053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4596.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4597 (.I0(\XII[18][3] ), .I1(\XII[19][3] ), .I2(n51770), 
            .O(n3054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4597.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4598 (.I0(n3054), .I1(n3053), .I2(n2959), .I3(n2953), 
            .O(n3055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4598.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4599 (.I0(n3055), .I1(n3052), .I2(n2967), .I3(n2966), 
            .O(n3056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__4599.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__4600 (.I0(n3049), .I1(n2959), .I2(n2967), .I3(n3056), 
            .O(n3057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd700 */ ;
    defparam LUT__4600.LUTMASK = 16'hd700;
    EFX_LUT4 LUT__4601 (.I0(n3043), .I1(n3057), .O(n3058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__4601.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__4602 (.I0(n2983), .I1(\PC[3] ), .I2(n2967), .I3(n2989), 
            .O(n3059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__4602.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__4603 (.I0(n3059), .I1(n2980), .I2(n2986), .O(n3060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__4603.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__4604 (.I0(\PC[3] ), .I1(n51758), .I2(n51838), .I3(n2981), 
            .O(n3061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4604.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4605 (.I0(n3061), .I1(n2986), .O(n3062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4605.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4606 (.I0(n3043), .I1(n2981), .I2(n3057), .I3(n3062), 
            .O(n3063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__4606.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__4607 (.I0(n2985), .I1(n3058), .I2(n3060), .I3(n3063), 
            .O(n523_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__4607.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__4608 (.I0(\XII[31][2] ), .I1(\XII[29][2] ), .I2(n2954), 
            .I3(n2953), .O(n3064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4608.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4609 (.I0(\XII[28][2] ), .I1(\XII[30][2] ), .I2(n2954), 
            .I3(n3064), .O(n3065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4609.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4610 (.I0(\XII[27][2] ), .I1(\XII[25][2] ), .I2(n2954), 
            .I3(n2953), .O(n3066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4610.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4611 (.I0(\XII[26][2] ), .I1(\XII[24][2] ), .I2(n2954), 
            .I3(n3066), .O(n3067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4611.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4612 (.I0(n3067), .I1(n3065), .I2(n2959), .I3(n2967), 
            .O(n3068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4612.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4613 (.I0(\XII[15][2] ), .I1(\XII[14][2] ), .I2(n2954), 
            .I3(n2953), .O(n3069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4613.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4614 (.I0(\XII[13][2] ), .I1(\XII[12][2] ), .I2(n2953), 
            .I3(n2954), .O(n3070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4614.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4615 (.I0(n3069), .I1(n3070), .I2(n2959), .O(n3071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4615.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4616 (.I0(\XII[9][2] ), .I1(\XII[8][2] ), .I2(n2954), 
            .O(n3072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4616.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4617 (.I0(\XII[11][2] ), .I1(\XII[10][2] ), .I2(n2954), 
            .O(n3073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4617.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4618 (.I0(n3073), .I1(n3072), .I2(n2959), .I3(n2953), 
            .O(n3074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4618.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4619 (.I0(\XII[5][2] ), .I1(\XII[4][2] ), .I2(n2953), 
            .I3(n2954), .O(n3075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4619.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4620 (.I0(\XII[7][2] ), .I1(\XII[6][2] ), .I2(n2954), 
            .I3(n2953), .O(n3076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4620.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4621 (.I0(\XII[1][2] ), .I1(\XII[0][2] ), .I2(STAGE2_EN), 
            .I3(n51770), .O(n3077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333 */ ;
    defparam LUT__4621.LUTMASK = 16'h5333;
    EFX_LUT4 LUT__4622 (.I0(\XII[2][2] ), .I1(\XII[3][2] ), .I2(n51770), 
            .O(n3078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4622.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4623 (.I0(n3078), .I1(n3077), .I2(n2953), .O(n3079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__4623.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__4624 (.I0(n3076), .I1(n3075), .I2(n3079), .I3(n2959), 
            .O(n3080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4624.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4625 (.I0(n3074), .I1(n3071), .I2(n3080), .I3(n2967), 
            .O(n3081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4625.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4626 (.I0(\XII[19][2] ), .I1(\XII[17][2] ), .I2(n2954), 
            .I3(n2953), .O(n3082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4626.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4627 (.I0(\XII[16][2] ), .I1(\XII[18][2] ), .I2(n2954), 
            .I3(n3082), .O(n3083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4627.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4628 (.I0(\XII[23][2] ), .I1(\XII[21][2] ), .I2(n2954), 
            .I3(n2953), .O(n3084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4628.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4629 (.I0(\XII[22][2] ), .I1(\XII[20][2] ), .I2(n2954), 
            .I3(n3084), .O(n3085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4629.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4630 (.I0(n3085), .I1(n3083), .I2(n2967), .I3(n2959), 
            .O(n3086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4630.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4631 (.I0(n3068), .I1(n3086), .I2(n3081), .I3(n2966), 
            .O(n3087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4631.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4632 (.I0(\PC[2] ), .I1(n51762), .I2(n51838), .I3(n2986), 
            .O(n3088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4632.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4633 (.I0(n2983), .I1(\PC[2] ), .I2(n2959), .I3(n2989), 
            .O(n3089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__4633.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__4634 (.I0(n2980), .I1(n2986), .O(n3090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__4634.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__4635 (.I0(n3089), .I1(n3090), .I2(n2981), .I3(n3088), 
            .O(n3091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4635.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4636 (.I0(n3087), .I1(n2987), .I2(n3091), .O(n524_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__4636.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__4637 (.I0(\XII[31][5] ), .I1(\XII[29][5] ), .I2(n2954), 
            .I3(n2953), .O(n3092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4637.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4638 (.I0(\XII[28][5] ), .I1(\XII[30][5] ), .I2(n2954), 
            .I3(n3092), .O(n3093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4638.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4639 (.I0(\XII[27][5] ), .I1(\XII[25][5] ), .I2(n2954), 
            .I3(n2953), .O(n3094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4639.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4640 (.I0(\XII[26][5] ), .I1(\XII[24][5] ), .I2(n2954), 
            .I3(n3094), .O(n3095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4640.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4641 (.I0(n3095), .I1(n3093), .I2(n2959), .I3(n2967), 
            .O(n3096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4641.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4642 (.I0(\XII[15][5] ), .I1(\XII[14][5] ), .I2(n2954), 
            .I3(n2953), .O(n3097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4642.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4643 (.I0(\XII[13][5] ), .I1(\XII[12][5] ), .I2(n2953), 
            .I3(n2954), .O(n3098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4643.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4644 (.I0(n3097), .I1(n3098), .I2(n2959), .O(n3099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4644.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4645 (.I0(\XII[9][5] ), .I1(\XII[8][5] ), .I2(n2954), 
            .O(n3100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4645.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4646 (.I0(\XII[11][5] ), .I1(\XII[10][5] ), .I2(n2954), 
            .O(n3101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4646.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4647 (.I0(n3101), .I1(n3100), .I2(n2959), .I3(n2953), 
            .O(n3102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4647.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4648 (.I0(\XII[5][5] ), .I1(\XII[4][5] ), .I2(n2953), 
            .I3(n2954), .O(n3103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4648.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4649 (.I0(\XII[7][5] ), .I1(\XII[6][5] ), .I2(n2954), 
            .I3(n2953), .O(n3104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4649.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4653 (.I0(n3104), .I1(n3103), .I2(n3107), .I3(n2959), 
            .O(n3108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4653.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4654 (.I0(n3102), .I1(n3099), .I2(n3108), .I3(n2967), 
            .O(n3109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4654.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4655 (.I0(\XII[19][5] ), .I1(\XII[17][5] ), .I2(n2954), 
            .I3(n2953), .O(n3110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4655.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4656 (.I0(\XII[16][5] ), .I1(\XII[18][5] ), .I2(n2954), 
            .I3(n3110), .O(n3111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4656.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4657 (.I0(\XII[23][5] ), .I1(\XII[21][5] ), .I2(n2954), 
            .I3(n2953), .O(n3112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4657.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4658 (.I0(\XII[22][5] ), .I1(\XII[20][5] ), .I2(n2954), 
            .I3(n3112), .O(n3113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4658.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4659 (.I0(n3113), .I1(n3111), .I2(n2967), .I3(n2959), 
            .O(n3114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4659.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4660 (.I0(n3096), .I1(n3114), .I2(n3109), .I3(n2966), 
            .O(n3115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4660.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4661 (.I0(\PC[5] ), .I1(n51750), .I2(n51838), .I3(n2986), 
            .O(n3116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4661.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4662 (.I0(\PC[5] ), .I1(n51834), .I2(n51750), .I3(n51842), 
            .O(n3117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__4662.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__4663 (.I0(n2980), .I1(STAGE2_EN), .O(n3118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4663.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4664 (.I0(n3117), .I1(n51838), .I2(n3118), .O(n3119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__4664.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__4665 (.I0(n2983), .I1(n2980), .I2(n2986), .O(n3120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__4665.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__4666 (.I0(n3119), .I1(n3120), .I2(n2981), .I3(n3116), 
            .O(n3121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4666.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4667 (.I0(n3115), .I1(n2987), .I2(n3121), .O(n521_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__4667.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__4668 (.I0(\XII[31][1] ), .I1(\XII[29][1] ), .I2(n2954), 
            .I3(n2953), .O(n3122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4668.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4669 (.I0(\XII[28][1] ), .I1(\XII[30][1] ), .I2(n2954), 
            .I3(n3122), .O(n3123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4669.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4670 (.I0(\XII[27][1] ), .I1(\XII[25][1] ), .I2(n2954), 
            .I3(n2953), .O(n3124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4670.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4671 (.I0(\XII[26][1] ), .I1(\XII[24][1] ), .I2(n2954), 
            .I3(n3124), .O(n3125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4671.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4672 (.I0(n3125), .I1(n3123), .I2(n2959), .I3(n2967), 
            .O(n3126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4672.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4673 (.I0(\XII[15][1] ), .I1(\XII[14][1] ), .I2(n2954), 
            .I3(n2953), .O(n3127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4673.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4674 (.I0(\XII[13][1] ), .I1(\XII[12][1] ), .I2(n2953), 
            .I3(n2954), .O(n3128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4674.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4675 (.I0(n3127), .I1(n3128), .I2(n2959), .O(n3129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4675.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4676 (.I0(\XII[9][1] ), .I1(\XII[8][1] ), .I2(n2954), 
            .O(n3130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4676.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4677 (.I0(\XII[11][1] ), .I1(\XII[10][1] ), .I2(n2954), 
            .O(n3131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4677.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4678 (.I0(n3131), .I1(n3130), .I2(n2959), .I3(n2953), 
            .O(n3132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4678.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4679 (.I0(\XII[5][1] ), .I1(\XII[4][1] ), .I2(n2953), 
            .I3(n2954), .O(n3133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4679.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4680 (.I0(\XII[7][1] ), .I1(\XII[6][1] ), .I2(n2954), 
            .I3(n2953), .O(n3134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4680.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4681 (.I0(\XII[1][1] ), .I1(\XII[0][1] ), .I2(STAGE2_EN), 
            .I3(n51770), .O(n3135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333 */ ;
    defparam LUT__4681.LUTMASK = 16'h5333;
    EFX_LUT4 LUT__4682 (.I0(\XII[2][1] ), .I1(\XII[3][1] ), .I2(n51770), 
            .O(n3136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4682.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4683 (.I0(n3136), .I1(n3135), .I2(n2953), .O(n3137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__4683.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__4684 (.I0(n3134), .I1(n3133), .I2(n3137), .I3(n2959), 
            .O(n3138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4684.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4685 (.I0(n3132), .I1(n3129), .I2(n3138), .I3(n2967), 
            .O(n3139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4685.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4686 (.I0(\XII[19][1] ), .I1(\XII[17][1] ), .I2(n2954), 
            .I3(n2953), .O(n3140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4686.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4687 (.I0(\XII[16][1] ), .I1(\XII[18][1] ), .I2(n2954), 
            .I3(n3140), .O(n3141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4687.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4688 (.I0(\XII[23][1] ), .I1(\XII[21][1] ), .I2(n2954), 
            .I3(n2953), .O(n3142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4688.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4689 (.I0(\XII[22][1] ), .I1(\XII[20][1] ), .I2(n2954), 
            .I3(n3142), .O(n3143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4689.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4690 (.I0(n3143), .I1(n3141), .I2(n2967), .I3(n2959), 
            .O(n3144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4690.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4691 (.I0(n3126), .I1(n3144), .I2(n3139), .I3(n2966), 
            .O(n3145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4691.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4692 (.I0(\PC[1] ), .I1(n51766), .I2(n51838), .I3(n2986), 
            .O(n3146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4692.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4693 (.I0(n2983), .I1(\PC[1] ), .I2(n2953), .I3(n2989), 
            .O(n3147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__4693.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__4694 (.I0(n3147), .I1(n3090), .I2(n2981), .I3(n3146), 
            .O(n3148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4694.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4695 (.I0(n3145), .I1(n2987), .I2(n3148), .O(n525_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__4695.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__4696 (.I0(STAGE2_EN), .I1(n51790), .O(\INSTRUCTION[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4696.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4697 (.I0(STAGE2_EN), .I1(n51786), .O(\INSTRUCTION[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4697.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4698 (.I0(\XII[15][0] ), .I1(\XII[13][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4698.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4699 (.I0(\XII[14][0] ), .I1(\XII[12][0] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4699.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4700 (.I0(STAGE2_EN), .I1(n51782), .O(\INSTRUCTION[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4700.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4701 (.I0(\XII[11][0] ), .I1(\XII[9][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4701.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4702 (.I0(\XII[10][0] ), .I1(\XII[8][0] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4702.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4703 (.I0(STAGE2_EN), .I1(n51778), .O(\INSTRUCTION[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4703.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4704 (.I0(\INSTRUCTION[17] ), .I1(n3152), .I2(n3151), 
            .I3(\INSTRUCTION[18] ), .O(n3153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__4704.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__4705 (.I0(n3150), .I1(n3149), .I2(\INSTRUCTION[17] ), 
            .I3(n3153), .O(n3154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__4705.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__4706 (.I0(STAGE2_EN), .I1(n51774), .O(\INSTRUCTION[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4706.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4707 (.I0(n2986), .I1(n3026), .I2(n51842), .O(n3155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4707.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4708 (.I0(\INSTRUCTION[19] ), .I1(n3154), .I2(n51766), 
            .I3(n3155), .O(n3156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__4708.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__4709 (.I0(\XII[31][0] ), .I1(\XII[29][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4709.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4710 (.I0(\XII[30][0] ), .I1(\XII[28][0] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4710.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4711 (.I0(\XII[27][0] ), .I1(\XII[25][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4711.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4712 (.I0(\XII[26][0] ), .I1(\XII[24][0] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4712.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4713 (.I0(\INSTRUCTION[17] ), .I1(n3160), .I2(n3159), 
            .I3(\INSTRUCTION[18] ), .O(n3161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__4713.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__4714 (.I0(n3158), .I1(n3157), .I2(\INSTRUCTION[17] ), 
            .I3(n3161), .O(n3162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__4714.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__4715 (.I0(\XII[7][0] ), .I1(\XII[3][0] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n3163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4715.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4716 (.I0(\XII[5][0] ), .I1(\XII[1][0] ), .I2(n51786), 
            .I3(n3163), .O(n3164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4716.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4717 (.I0(\XII[6][0] ), .I1(\XII[2][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n3165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4717.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4718 (.I0(\XII[4][0] ), .I1(\XII[0][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(n3165), .O(n3166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4718.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4719 (.I0(n3166), .I1(n3164), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n3167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__4719.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__4720 (.I0(\XII[23][0] ), .I1(\XII[19][0] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n3168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4720.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4721 (.I0(\XII[21][0] ), .I1(\XII[17][0] ), .I2(n51786), 
            .I3(n3168), .O(n3169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4721.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4722 (.I0(\XII[22][0] ), .I1(\XII[18][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n3170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4722.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4723 (.I0(\XII[20][0] ), .I1(\XII[16][0] ), .I2(\INSTRUCTION[16] ), 
            .I3(n3170), .O(n3171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4723.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4724 (.I0(n3171), .I1(n3169), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n3172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__4724.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__4725 (.I0(n3162), .I1(n3172), .I2(n3167), .I3(\INSTRUCTION[19] ), 
            .O(n3173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4725.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4726 (.I0(n51826), .I1(n2983), .O(n3174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4726.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4727 (.I0(n3155), .I1(n3173), .I2(n3174), .I3(n3156), 
            .O(n574_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__4727.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__4728 (.I0(\XII[31][0] ), .I1(\XII[29][0] ), .I2(n2954), 
            .I3(n2953), .O(n3175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4728.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4729 (.I0(\XII[28][0] ), .I1(\XII[30][0] ), .I2(n2954), 
            .I3(n3175), .O(n3176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4729.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4730 (.I0(\XII[27][0] ), .I1(\XII[25][0] ), .I2(n2954), 
            .I3(n2953), .O(n3177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4730.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4731 (.I0(\XII[26][0] ), .I1(\XII[24][0] ), .I2(n2954), 
            .I3(n3177), .O(n3178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4731.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4732 (.I0(n3178), .I1(n3176), .I2(n2959), .I3(n2967), 
            .O(n3179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4732.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4733 (.I0(\XII[15][0] ), .I1(\XII[14][0] ), .I2(n2954), 
            .I3(n2953), .O(n3180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4733.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4734 (.I0(\XII[13][0] ), .I1(\XII[12][0] ), .I2(n2953), 
            .I3(n2954), .O(n3181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4734.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4735 (.I0(n3180), .I1(n3181), .I2(n2959), .O(n3182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4735.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4736 (.I0(\XII[9][0] ), .I1(\XII[8][0] ), .I2(n2954), 
            .O(n3183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4736.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4737 (.I0(\XII[11][0] ), .I1(\XII[10][0] ), .I2(n2954), 
            .O(n3184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4737.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4738 (.I0(n3184), .I1(n3183), .I2(n2959), .I3(n2953), 
            .O(n3185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4738.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4739 (.I0(\XII[5][0] ), .I1(\XII[4][0] ), .I2(n2953), 
            .I3(n2954), .O(n3186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4739.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4740 (.I0(\XII[7][0] ), .I1(\XII[6][0] ), .I2(n2954), 
            .I3(n2953), .O(n3187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4740.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4741 (.I0(\XII[1][0] ), .I1(\XII[0][0] ), .I2(STAGE2_EN), 
            .I3(n51770), .O(n3188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333 */ ;
    defparam LUT__4741.LUTMASK = 16'h5333;
    EFX_LUT4 LUT__4742 (.I0(\XII[2][0] ), .I1(\XII[3][0] ), .I2(n51770), 
            .O(n3189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4742.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4743 (.I0(n3189), .I1(n3188), .I2(n2953), .O(n3190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__4743.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__4744 (.I0(n3187), .I1(n3186), .I2(n3190), .I3(n2959), 
            .O(n3191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4744.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4745 (.I0(n3185), .I1(n3182), .I2(n3191), .I3(n2967), 
            .O(n3192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4745.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4746 (.I0(\XII[19][0] ), .I1(\XII[17][0] ), .I2(n2954), 
            .I3(n2953), .O(n3193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4746.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4747 (.I0(\XII[16][0] ), .I1(\XII[18][0] ), .I2(n2954), 
            .I3(n3193), .O(n3194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4747.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4748 (.I0(\XII[23][0] ), .I1(\XII[21][0] ), .I2(n2954), 
            .I3(n2953), .O(n3195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4748.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4749 (.I0(\XII[22][0] ), .I1(\XII[20][0] ), .I2(n2954), 
            .I3(n3195), .O(n3196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4749.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4750 (.I0(n3196), .I1(n3194), .I2(n2967), .I3(n2959), 
            .O(n3197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4750.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4751 (.I0(n3179), .I1(n3197), .I2(n3192), .I3(n2966), 
            .O(n3198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4751.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4752 (.I0(\PC[0] ), .I1(n51770), .I2(n51838), .I3(n2986), 
            .O(n3199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__4752.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__4753 (.I0(\PC[0] ), .I1(n2983), .I2(n2954), .I3(n2989), 
            .O(n3200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4753.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4754 (.I0(n3200), .I1(n3090), .I2(n2981), .I3(n3199), 
            .O(n3201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4754.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4755 (.I0(n3198), .I1(n2987), .I2(n3201), .O(n526_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__4755.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__4756 (.I0(n2989), .I1(n51826), .I2(STAGE2_EN), .O(n3202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__4756.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__4757 (.I0(n3202), .I1(n51830), .I2(n2982), .O(n3203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4757.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4758 (.I0(n3198), .I1(n2954), .I2(n3203), .O(n541_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__4758.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__4759 (.I0(n51730), .I1(n51794), .I2(n51802), .I3(n51798), 
            .O(n3204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fb3 */ ;
    defparam LUT__4759.LUTMASK = 16'h0fb3;
    EFX_LUT4 LUT__4760 (.I0(n51798), .I1(n51802), .I2(n51730), .I3(n51834), 
            .O(n3205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__4760.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__4761 (.I0(n3205), .I1(n51830), .I2(STAGE2_EN), .O(n3206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4761.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4762 (.I0(n3204), .I1(n2982), .I2(n3206), .I3(n3202), 
            .O(n531_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__4762.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__4763 (.I0(n51830), .I1(n51794), .I2(\DATA_FORMAT[0] ), 
            .I3(n51798), .O(n3207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__4763.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__4764 (.I0(n3207), .I1(STAGE2_EN), .I2(n51802), .O(n49404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4764.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4765 (.I0(n51834), .I1(n51794), .I2(n2989), .O(n3208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4765.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4766 (.I0(n51794), .I1(n51798), .I2(n51834), .O(n3209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__4766.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__4767 (.I0(n2989), .I1(n3209), .I2(n51830), .I3(STAGE2_EN), 
            .O(n3210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__4767.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__4768 (.I0(n3210), .I1(n2986), .I2(n30664), .O(n3211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4768.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4769 (.I0(n3208), .I1(STAGE2_EN), .I2(n51830), .I3(n3211), 
            .O(ceg_net35296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff */ ;
    defparam LUT__4769.LUTMASK = 16'h40ff;
    EFX_LUT4 LUT__4770 (.I0(STAGE2_EN), .I1(n51822), .O(\INSTRUCTION[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4770.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4771 (.I0(n3202), .I1(n3028), .I2(n30664), .O(n50065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__4771.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__4772 (.I0(\XII[31][6] ), .I1(\XII[29][6] ), .I2(n2954), 
            .I3(n2953), .O(n3212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4772.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4773 (.I0(\XII[28][6] ), .I1(\XII[30][6] ), .I2(n2954), 
            .I3(n3212), .O(n3213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4773.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4774 (.I0(\XII[27][6] ), .I1(\XII[25][6] ), .I2(n2954), 
            .I3(n2953), .O(n3214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4774.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4775 (.I0(\XII[26][6] ), .I1(\XII[24][6] ), .I2(n2954), 
            .I3(n3214), .O(n3215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4775.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4776 (.I0(n3215), .I1(n3213), .I2(n2959), .I3(n2967), 
            .O(n3216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4776.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4777 (.I0(\XII[15][6] ), .I1(\XII[14][6] ), .I2(n2954), 
            .I3(n2953), .O(n3217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4777.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4778 (.I0(\XII[13][6] ), .I1(\XII[12][6] ), .I2(n2953), 
            .I3(n2954), .O(n3218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4778.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4779 (.I0(n3217), .I1(n3218), .I2(n2959), .O(n3219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4779.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4780 (.I0(\XII[9][6] ), .I1(\XII[8][6] ), .I2(n2954), 
            .O(n3220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4780.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4781 (.I0(\XII[11][6] ), .I1(\XII[10][6] ), .I2(n2954), 
            .O(n3221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4781.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4782 (.I0(n3221), .I1(n3220), .I2(n2959), .I3(n2953), 
            .O(n3222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4782.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4783 (.I0(\XII[5][6] ), .I1(\XII[4][6] ), .I2(n2953), 
            .I3(n2954), .O(n3223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4783.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4784 (.I0(\XII[7][6] ), .I1(\XII[6][6] ), .I2(n2954), 
            .I3(n2953), .O(n3224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4784.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4788 (.I0(n3224), .I1(n3223), .I2(n3227), .I3(n2959), 
            .O(n3228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4788.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4789 (.I0(n3222), .I1(n3219), .I2(n3228), .I3(n2967), 
            .O(n3229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4789.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4790 (.I0(\XII[19][6] ), .I1(\XII[17][6] ), .I2(n2954), 
            .I3(n2953), .O(n3230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4790.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4791 (.I0(\XII[16][6] ), .I1(\XII[18][6] ), .I2(n2954), 
            .I3(n3230), .O(n3231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4791.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4792 (.I0(\XII[23][6] ), .I1(\XII[21][6] ), .I2(n2954), 
            .I3(n2953), .O(n3232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4792.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4793 (.I0(\XII[22][6] ), .I1(\XII[20][6] ), .I2(n2954), 
            .I3(n3232), .O(n3233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4793.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4794 (.I0(n3233), .I1(n3231), .I2(n2967), .I3(n2959), 
            .O(n3234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4794.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4795 (.I0(n3216), .I1(n3234), .I2(n3229), .I3(n2966), 
            .O(n3235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4795.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4796 (.I0(\PC[6] ), .I1(n51746), .I2(n51838), .I3(n2986), 
            .O(n3236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4796.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4797 (.I0(\PC[6] ), .I1(n51834), .I2(n51746), .I3(n51842), 
            .O(n3237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__4797.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__4798 (.I0(n3237), .I1(n51838), .I2(n3118), .O(n3238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__4798.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__4799 (.I0(n3238), .I1(n3120), .I2(n2981), .I3(n3236), 
            .O(n3239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4799.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4800 (.I0(n3235), .I1(n2987), .I2(n3239), .O(n520_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__4800.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__4801 (.I0(\XII[31][7] ), .I1(\XII[29][7] ), .I2(n2954), 
            .I3(n2953), .O(n3240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4801.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4802 (.I0(\XII[28][7] ), .I1(\XII[30][7] ), .I2(n2954), 
            .I3(n3240), .O(n3241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4802.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4803 (.I0(\XII[27][7] ), .I1(\XII[25][7] ), .I2(n2954), 
            .I3(n2953), .O(n3242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4803.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4804 (.I0(\XII[26][7] ), .I1(\XII[24][7] ), .I2(n2954), 
            .I3(n3242), .O(n3243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4804.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4805 (.I0(n3243), .I1(n3241), .I2(n2959), .I3(n2967), 
            .O(n3244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4805.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4806 (.I0(\XII[15][7] ), .I1(\XII[14][7] ), .I2(n2954), 
            .I3(n2953), .O(n3245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4806.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4807 (.I0(\XII[13][7] ), .I1(\XII[12][7] ), .I2(n2953), 
            .I3(n2954), .O(n3246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4807.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4808 (.I0(n3245), .I1(n3246), .I2(n2959), .O(n3247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4808.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4809 (.I0(\XII[9][7] ), .I1(\XII[8][7] ), .I2(n2954), 
            .O(n3248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4809.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4810 (.I0(\XII[11][7] ), .I1(\XII[10][7] ), .I2(n2954), 
            .O(n3249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4810.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4811 (.I0(n3249), .I1(n3248), .I2(n2959), .I3(n2953), 
            .O(n3250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4811.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4812 (.I0(\XII[5][7] ), .I1(\XII[4][7] ), .I2(n2953), 
            .I3(n2954), .O(n3251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4812.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4813 (.I0(\XII[7][7] ), .I1(\XII[6][7] ), .I2(n2954), 
            .I3(n2953), .O(n3252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4813.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4817 (.I0(n3252), .I1(n3251), .I2(n3255), .I3(n2959), 
            .O(n3256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4817.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4818 (.I0(n3250), .I1(n3247), .I2(n3256), .I3(n2967), 
            .O(n3257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4818.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4819 (.I0(\XII[19][7] ), .I1(\XII[17][7] ), .I2(n2954), 
            .I3(n2953), .O(n3258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4819.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4820 (.I0(\XII[16][7] ), .I1(\XII[18][7] ), .I2(n2954), 
            .I3(n3258), .O(n3259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4820.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4821 (.I0(\XII[23][7] ), .I1(\XII[21][7] ), .I2(n2954), 
            .I3(n2953), .O(n3260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4821.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4822 (.I0(\XII[22][7] ), .I1(\XII[20][7] ), .I2(n2954), 
            .I3(n3260), .O(n3261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4822.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4823 (.I0(n3261), .I1(n3259), .I2(n2967), .I3(n2959), 
            .O(n3262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4823.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4824 (.I0(n3244), .I1(n3262), .I2(n3257), .I3(n2966), 
            .O(n3263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4824.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4825 (.I0(\PC[7] ), .I1(n51742), .I2(n51838), .I3(n2986), 
            .O(n3264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4825.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4826 (.I0(\PC[7] ), .I1(n51834), .I2(n51742), .I3(n51842), 
            .O(n3265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__4826.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__4827 (.I0(n3265), .I1(n51838), .I2(n3118), .O(n3266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__4827.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__4828 (.I0(n3266), .I1(n3120), .I2(n2981), .I3(n3264), 
            .O(n3267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4828.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4829 (.I0(n3263), .I1(n2987), .I2(n3267), .O(n519_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__4829.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__4830 (.I0(\XI[31][8] ), .I1(\XI[29][8] ), .I2(n2954), 
            .I3(n2953), .O(n3268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4830.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4831 (.I0(\XI[28][8] ), .I1(\XI[30][8] ), .I2(n2954), 
            .I3(n3268), .O(n3269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4831.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4832 (.I0(\XI[27][8] ), .I1(\XI[25][8] ), .I2(n2954), 
            .I3(n2953), .O(n3270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4832.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4833 (.I0(\XI[26][8] ), .I1(\XI[24][8] ), .I2(n2954), 
            .I3(n3270), .O(n3271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4833.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4834 (.I0(n3271), .I1(n3269), .I2(n2959), .I3(n2967), 
            .O(n3272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4834.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4835 (.I0(\XI[15][8] ), .I1(\XI[14][8] ), .I2(n2954), 
            .I3(n2953), .O(n3273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4835.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4836 (.I0(\XI[13][8] ), .I1(\XI[12][8] ), .I2(n2953), 
            .I3(n2954), .O(n3274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4836.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4837 (.I0(n3273), .I1(n3274), .I2(n2959), .O(n3275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4837.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4838 (.I0(\XI[9][8] ), .I1(\XI[8][8] ), .I2(n2954), 
            .O(n3276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4838.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4839 (.I0(\XI[11][8] ), .I1(\XI[10][8] ), .I2(n2954), 
            .O(n3277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4839.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4840 (.I0(n3277), .I1(n3276), .I2(n2959), .I3(n2953), 
            .O(n3278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4840.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4841 (.I0(\XI[5][8] ), .I1(\XI[4][8] ), .I2(n2953), 
            .I3(n2954), .O(n3279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4841.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4842 (.I0(\XI[7][8] ), .I1(\XI[6][8] ), .I2(n2954), 
            .I3(n2953), .O(n3280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4842.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4846 (.I0(n3280), .I1(n3279), .I2(n3283), .I3(n2959), 
            .O(n3284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4846.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4847 (.I0(n3278), .I1(n3275), .I2(n3284), .I3(n2967), 
            .O(n3285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4847.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4848 (.I0(\XI[19][8] ), .I1(\XI[17][8] ), .I2(n2954), 
            .I3(n2953), .O(n3286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4848.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4849 (.I0(\XI[16][8] ), .I1(\XI[18][8] ), .I2(n2954), 
            .I3(n3286), .O(n3287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4849.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4850 (.I0(\XI[23][8] ), .I1(\XI[21][8] ), .I2(n2954), 
            .I3(n2953), .O(n3288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4850.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4851 (.I0(\XI[22][8] ), .I1(\XI[20][8] ), .I2(n2954), 
            .I3(n3288), .O(n3289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4851.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4852 (.I0(n3289), .I1(n3287), .I2(n2967), .I3(n2959), 
            .O(n3290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4852.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4853 (.I0(n3272), .I1(n3290), .I2(n3285), .I3(n2966), 
            .O(n3291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4853.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4854 (.I0(\PC[8] ), .I1(n51738), .I2(n51838), .I3(n2986), 
            .O(n3292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4854.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4855 (.I0(\PC[8] ), .I1(n51834), .I2(n51738), .I3(n51842), 
            .O(n3293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__4855.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__4856 (.I0(n3293), .I1(n51838), .I2(n3118), .O(n3294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__4856.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__4857 (.I0(n3294), .I1(n3120), .I2(n2981), .I3(n3292), 
            .O(n3295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4857.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4858 (.I0(n3291), .I1(n2987), .I2(n3295), .O(n518_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__4858.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__4859 (.I0(\PC[9] ), .I1(n51734), .I2(n51842), .O(n3296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4859.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4860 (.I0(n3296), .I1(n3118), .O(n3297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4860.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4861 (.I0(\XI[31][9] ), .I1(\XI[29][9] ), .I2(n2954), 
            .I3(n2953), .O(n3298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4861.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4862 (.I0(\XI[28][9] ), .I1(\XI[30][9] ), .I2(n2954), 
            .I3(n3298), .O(n3299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4862.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4863 (.I0(\XI[27][9] ), .I1(\XI[25][9] ), .I2(n2954), 
            .I3(n2953), .O(n3300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4863.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4864 (.I0(\XI[26][9] ), .I1(\XI[24][9] ), .I2(n2954), 
            .I3(n3300), .O(n3301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4864.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4865 (.I0(n3301), .I1(n3299), .I2(n2959), .I3(n2967), 
            .O(n3302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4865.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4866 (.I0(\XI[15][9] ), .I1(\XI[14][9] ), .I2(n2954), 
            .I3(n2953), .O(n3303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4866.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4867 (.I0(\XI[13][9] ), .I1(\XI[12][9] ), .I2(n2953), 
            .I3(n2954), .O(n3304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4867.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4868 (.I0(n3303), .I1(n3304), .I2(n2959), .O(n3305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4868.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4869 (.I0(\XI[9][9] ), .I1(\XI[8][9] ), .I2(n2954), 
            .O(n3306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4869.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4870 (.I0(\XI[11][9] ), .I1(\XI[10][9] ), .I2(n2954), 
            .O(n3307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4870.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4871 (.I0(n3307), .I1(n3306), .I2(n2959), .I3(n2953), 
            .O(n3308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4871.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4872 (.I0(\XI[5][9] ), .I1(\XI[4][9] ), .I2(n2953), 
            .I3(n2954), .O(n3309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4872.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4873 (.I0(\XI[7][9] ), .I1(\XI[6][9] ), .I2(n2954), 
            .I3(n2953), .O(n3310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4873.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4877 (.I0(n3310), .I1(n3309), .I2(n3313), .I3(n2959), 
            .O(n3314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4877.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4878 (.I0(n3308), .I1(n3305), .I2(n3314), .I3(n2967), 
            .O(n3315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4878.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4879 (.I0(\XI[19][9] ), .I1(\XI[17][9] ), .I2(n2954), 
            .I3(n2953), .O(n3316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4879.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4880 (.I0(\XI[16][9] ), .I1(\XI[18][9] ), .I2(n2954), 
            .I3(n3316), .O(n3317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4880.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4881 (.I0(\XI[23][9] ), .I1(\XI[21][9] ), .I2(n2954), 
            .I3(n2953), .O(n3318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4881.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4882 (.I0(\XI[22][9] ), .I1(\XI[20][9] ), .I2(n2954), 
            .I3(n3318), .O(n3319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4882.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4883 (.I0(n3319), .I1(n3317), .I2(n2967), .I3(n2959), 
            .O(n3320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4883.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4884 (.I0(n3302), .I1(n3320), .I2(n3315), .I3(n2966), 
            .O(n3321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4884.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4885 (.I0(\PC[9] ), .I1(n51734), .I2(n51838), .I3(n2981), 
            .O(n3322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4885.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4886 (.I0(n3322), .I1(n2986), .O(n3323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4886.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4887 (.I0(n3321), .I1(n3297), .I2(n3323), .I3(n2987), 
            .O(n517_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf5fc */ ;
    defparam LUT__4887.LUTMASK = 16'hf5fc;
    EFX_LUT4 LUT__4888 (.I0(\XI[31][10] ), .I1(\XI[29][10] ), .I2(n2954), 
            .I3(n2953), .O(n3324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4888.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4889 (.I0(\XI[28][10] ), .I1(\XI[30][10] ), .I2(n2954), 
            .I3(n3324), .O(n3325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4889.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4890 (.I0(\XI[27][10] ), .I1(\XI[25][10] ), .I2(n2954), 
            .I3(n2953), .O(n3326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4890.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4891 (.I0(\XI[26][10] ), .I1(\XI[24][10] ), .I2(n2954), 
            .I3(n3326), .O(n3327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4891.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4892 (.I0(n3327), .I1(n3325), .I2(n2959), .I3(n2967), 
            .O(n3328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__4892.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__4893 (.I0(\XI[15][10] ), .I1(\XI[14][10] ), .I2(n2954), 
            .I3(n2953), .O(n3329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4893.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4894 (.I0(\XI[13][10] ), .I1(\XI[12][10] ), .I2(n2953), 
            .I3(n2954), .O(n3330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4894.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4895 (.I0(n3329), .I1(n3330), .I2(n2959), .O(n3331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4895.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4896 (.I0(\XI[9][10] ), .I1(\XI[8][10] ), .I2(n2954), 
            .O(n3332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4896.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4897 (.I0(\XI[11][10] ), .I1(\XI[10][10] ), .I2(n2954), 
            .O(n3333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4897.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4898 (.I0(n3333), .I1(n3332), .I2(n2959), .I3(n2953), 
            .O(n3334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4898.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4899 (.I0(\XI[5][10] ), .I1(\XI[4][10] ), .I2(n2953), 
            .I3(n2954), .O(n3335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4899.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4900 (.I0(\XI[7][10] ), .I1(\XI[6][10] ), .I2(n2954), 
            .I3(n2953), .O(n3336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4900.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4904 (.I0(n3336), .I1(n3335), .I2(n3339), .I3(n2959), 
            .O(n3340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4904.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4905 (.I0(n3334), .I1(n3331), .I2(n3340), .I3(n2967), 
            .O(n3341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4905.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4906 (.I0(\XI[19][10] ), .I1(\XI[17][10] ), .I2(n2954), 
            .I3(n2953), .O(n3342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4906.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4907 (.I0(\XI[16][10] ), .I1(\XI[18][10] ), .I2(n2954), 
            .I3(n3342), .O(n3343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__4907.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__4908 (.I0(\XI[23][10] ), .I1(\XI[21][10] ), .I2(n2954), 
            .I3(n2953), .O(n3344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4908.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4909 (.I0(\XI[22][10] ), .I1(\XI[20][10] ), .I2(n2954), 
            .I3(n3344), .O(n3345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4909.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4910 (.I0(n3345), .I1(n3343), .I2(n2967), .I3(n2959), 
            .O(n3346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4910.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4911 (.I0(n3328), .I1(n3346), .I2(n3341), .I3(n2966), 
            .O(n3347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4911.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4912 (.I0(\PC[10] ), .I1(n51730), .I2(n51838), .I3(n2986), 
            .O(n3348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4912.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4913 (.I0(\PC[10] ), .I1(n51834), .I2(n51730), .I3(n51842), 
            .O(n3349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__4913.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__4914 (.I0(n3349), .I1(n51838), .I2(n3118), .O(n3350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__4914.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__4915 (.I0(n3350), .I1(n3120), .I2(n2981), .I3(n3348), 
            .O(n3351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__4915.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__4916 (.I0(n3347), .I1(n2987), .I2(n3351), .O(n516_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__4916.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__4917 (.I0(\XI[18][11] ), .I1(\XI[19][11] ), .I2(n51770), 
            .O(n3352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4917.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4918 (.I0(\XI[16][11] ), .I1(\XI[17][11] ), .I2(n51770), 
            .O(n3353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4918.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4919 (.I0(n3352), .I1(n3353), .I2(n2959), .I3(n2953), 
            .O(n3354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__4919.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__4920 (.I0(\XI[21][11] ), .I1(\XI[20][11] ), .I2(n2953), 
            .I3(n2954), .O(n3355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4920.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4921 (.I0(\XI[23][11] ), .I1(\XI[22][11] ), .I2(n51770), 
            .O(n3356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4921.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4922 (.I0(n3356), .I1(n3354), .I2(n3355), .I3(n2959), 
            .O(n3357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__4922.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__4923 (.I0(\XI[25][11] ), .I1(\XI[24][11] ), .I2(n2954), 
            .O(n3358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4923.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4924 (.I0(\XI[27][11] ), .I1(\XI[26][11] ), .I2(n2954), 
            .O(n3359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4924.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4925 (.I0(n3359), .I1(n3358), .I2(n2959), .I3(n2953), 
            .O(n3360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4925.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4926 (.I0(\XI[31][11] ), .I1(\XI[30][11] ), .I2(n2954), 
            .O(n3361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4926.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4927 (.I0(\XI[29][11] ), .I1(\XI[28][11] ), .I2(n2954), 
            .O(n3362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4927.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4928 (.I0(n3362), .I1(n3361), .I2(n2953), .I3(n2959), 
            .O(n3363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__4928.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__4929 (.I0(n3360), .I1(n3363), .I2(n3357), .I3(n2967), 
            .O(n3364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4929.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4930 (.I0(\XI[15][11] ), .I1(\XI[14][11] ), .I2(n2954), 
            .I3(n2953), .O(n3365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4930.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4931 (.I0(\XI[13][11] ), .I1(\XI[12][11] ), .I2(n2953), 
            .I3(n2954), .O(n3366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4931.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4932 (.I0(n3365), .I1(n3366), .I2(n2959), .O(n3367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4932.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4933 (.I0(\XI[9][11] ), .I1(\XI[8][11] ), .I2(n2954), 
            .O(n3368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4933.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4934 (.I0(\XI[11][11] ), .I1(\XI[10][11] ), .I2(n2954), 
            .O(n3369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4934.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4935 (.I0(n3369), .I1(n3368), .I2(n2959), .I3(n2953), 
            .O(n3370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4935.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4936 (.I0(\XI[5][11] ), .I1(\XI[4][11] ), .I2(n2953), 
            .I3(n2954), .O(n3371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4936.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4937 (.I0(\XI[7][11] ), .I1(\XI[6][11] ), .I2(n2954), 
            .I3(n2953), .O(n3372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4937.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4941 (.I0(n3372), .I1(n3371), .I2(n3375), .I3(n2959), 
            .O(n3376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4941.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4942 (.I0(n3370), .I1(n3367), .I2(n3376), .I3(n2967), 
            .O(n3377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4942.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4943 (.I0(n3377), .I1(n3364), .I2(n3029), .I3(n2966), 
            .O(n3378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__4943.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__4944 (.I0(n51726), .I1(n51838), .I2(n3029), .O(n3379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__4944.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__4945 (.I0(n51838), .I1(\PC[11] ), .I2(n3379), .I3(n2986), 
            .O(n3380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__4945.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__4946 (.I0(n3377), .I1(n3364), .I2(n2991), .I3(n2966), 
            .O(n3381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__4946.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__4947 (.I0(n2983), .I1(STAGE2_EN), .I2(n51830), .I3(n2990), 
            .O(n3382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__4947.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__4948 (.I0(n3382), .I1(n2986), .O(n3383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__4948.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__4949 (.I0(n2983), .I1(\PC[11] ), .I2(n3383), .O(n3384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__4949.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__4950 (.I0(n3381), .I1(n3384), .I2(n3378), .I3(n3380), 
            .O(n515_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__4950.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__4951 (.I0(\XI[18][12] ), .I1(\XI[19][12] ), .I2(n51770), 
            .O(n3385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4951.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4952 (.I0(\XI[16][12] ), .I1(\XI[17][12] ), .I2(n51770), 
            .O(n3386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4952.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4953 (.I0(n3385), .I1(n3386), .I2(n2959), .I3(n2953), 
            .O(n3387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__4953.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__4954 (.I0(\XI[21][12] ), .I1(\XI[20][12] ), .I2(n2953), 
            .I3(n2954), .O(n3388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4954.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4955 (.I0(\XI[23][12] ), .I1(\XI[22][12] ), .I2(n51770), 
            .O(n3389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4955.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4956 (.I0(n3389), .I1(n3387), .I2(n3388), .I3(n2959), 
            .O(n3390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__4956.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__4957 (.I0(\XI[25][12] ), .I1(\XI[24][12] ), .I2(n2954), 
            .O(n3391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4957.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4958 (.I0(\XI[27][12] ), .I1(\XI[26][12] ), .I2(n2954), 
            .O(n3392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4958.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4959 (.I0(n3392), .I1(n3391), .I2(n2959), .I3(n2953), 
            .O(n3393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4959.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4960 (.I0(\XI[31][12] ), .I1(\XI[30][12] ), .I2(n2954), 
            .O(n3394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4960.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4961 (.I0(\XI[29][12] ), .I1(\XI[28][12] ), .I2(n2954), 
            .O(n3395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4961.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4962 (.I0(n3395), .I1(n3394), .I2(n2953), .I3(n2959), 
            .O(n3396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__4962.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__4963 (.I0(n3393), .I1(n3396), .I2(n3390), .I3(n2967), 
            .O(n3397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4963.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4964 (.I0(\XI[15][12] ), .I1(\XI[14][12] ), .I2(n2954), 
            .I3(n2953), .O(n3398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4964.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4965 (.I0(\XI[13][12] ), .I1(\XI[12][12] ), .I2(n2953), 
            .I3(n2954), .O(n3399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4965.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4966 (.I0(n3398), .I1(n3399), .I2(n2959), .O(n3400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4966.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4967 (.I0(\XI[9][12] ), .I1(\XI[8][12] ), .I2(n2954), 
            .O(n3401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4967.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4968 (.I0(\XI[11][12] ), .I1(\XI[10][12] ), .I2(n2954), 
            .O(n3402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4968.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4969 (.I0(n3402), .I1(n3401), .I2(n2959), .I3(n2953), 
            .O(n3403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__4969.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__4970 (.I0(\XI[5][12] ), .I1(\XI[4][12] ), .I2(n2953), 
            .I3(n2954), .O(n3404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4970.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4971 (.I0(\XI[7][12] ), .I1(\XI[6][12] ), .I2(n2954), 
            .I3(n2953), .O(n3405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4971.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4975 (.I0(n3405), .I1(n3404), .I2(n3408), .I3(n2959), 
            .O(n3409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4975.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4976 (.I0(n3403), .I1(n3400), .I2(n3409), .I3(n2967), 
            .O(n3410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4976.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4977 (.I0(n3410), .I1(n3397), .I2(n3029), .I3(n2966), 
            .O(n3411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__4977.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__4978 (.I0(\PC[12] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__4978.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__4979 (.I0(n3410), .I1(n3397), .I2(n2991), .I3(n2966), 
            .O(n3413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__4979.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__4980 (.I0(n2983), .I1(\PC[12] ), .I2(n3383), .O(n3414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__4980.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__4981 (.I0(n3413), .I1(n3414), .I2(n3411), .I3(n3412), 
            .O(n514_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__4981.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__4982 (.I0(\XI[18][13] ), .I1(\XI[19][13] ), .I2(n51770), 
            .O(n3415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4982.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4983 (.I0(\XI[16][13] ), .I1(\XI[17][13] ), .I2(n51770), 
            .O(n3416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__4983.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__4984 (.I0(n3415), .I1(n3416), .I2(n2959), .I3(n2953), 
            .O(n3417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__4984.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__4985 (.I0(\XI[21][13] ), .I1(\XI[20][13] ), .I2(n2953), 
            .I3(n2954), .O(n3418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4985.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4986 (.I0(\XI[23][13] ), .I1(\XI[22][13] ), .I2(n51770), 
            .O(n3419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4986.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4987 (.I0(n3419), .I1(n3417), .I2(n3418), .I3(n2959), 
            .O(n3420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__4987.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__4988 (.I0(\XI[25][13] ), .I1(\XI[24][13] ), .I2(n2954), 
            .O(n3421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4988.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4989 (.I0(\XI[27][13] ), .I1(\XI[26][13] ), .I2(n2954), 
            .O(n3422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4989.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4990 (.I0(n3422), .I1(n3421), .I2(n2959), .I3(n2953), 
            .O(n3423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4990.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4991 (.I0(\XI[31][13] ), .I1(\XI[30][13] ), .I2(n2954), 
            .O(n3424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4991.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4992 (.I0(\XI[29][13] ), .I1(\XI[28][13] ), .I2(n2954), 
            .O(n3425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4992.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4993 (.I0(n3425), .I1(n3424), .I2(n2953), .I3(n2959), 
            .O(n3426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__4993.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__4994 (.I0(n3423), .I1(n3426), .I2(n3420), .I3(n2967), 
            .O(n3427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4994.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4995 (.I0(\XI[15][13] ), .I1(\XI[14][13] ), .I2(n2954), 
            .I3(n2953), .O(n3428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4995.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4996 (.I0(\XI[13][13] ), .I1(\XI[12][13] ), .I2(n2953), 
            .I3(n2954), .O(n3429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4996.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4997 (.I0(n3428), .I1(n3429), .I2(n2959), .O(n3430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4997.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4998 (.I0(\XI[9][13] ), .I1(\XI[8][13] ), .I2(n2954), 
            .O(n3431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4998.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4999 (.I0(\XI[11][13] ), .I1(\XI[10][13] ), .I2(n2954), 
            .O(n3432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4999.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5000 (.I0(n3432), .I1(n3431), .I2(n2959), .I3(n2953), 
            .O(n3433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5000.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5001 (.I0(\XI[5][13] ), .I1(\XI[4][13] ), .I2(n2953), 
            .I3(n2954), .O(n3434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5001.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5002 (.I0(\XI[7][13] ), .I1(\XI[6][13] ), .I2(n2954), 
            .I3(n2953), .O(n3435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5002.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5006 (.I0(n3435), .I1(n3434), .I2(n3438), .I3(n2959), 
            .O(n3439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5006.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5007 (.I0(n3433), .I1(n3430), .I2(n3439), .I3(n2967), 
            .O(n3440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5007.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5008 (.I0(n3440), .I1(n3427), .I2(n3029), .I3(n2966), 
            .O(n3441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5008.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5009 (.I0(\PC[13] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5009.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5010 (.I0(n3440), .I1(n3427), .I2(n2991), .I3(n2966), 
            .O(n3443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5010.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5011 (.I0(n2983), .I1(\PC[13] ), .I2(n3383), .O(n3444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5011.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5012 (.I0(n3443), .I1(n3444), .I2(n3441), .I3(n3442), 
            .O(n513_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5012.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5013 (.I0(\OPERATION[0] ), .I1(\OPERATION[1] ), .O(n3445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5013.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5014 (.I0(n3445), .I1(\OPERATION[3] ), .O(n1649_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5014.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5015 (.I0(STAGE3_EN), .I1(n221), .O(n30678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5015.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5016 (.I0(n1649_2), .I1(n30678), .O(n50476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__5016.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__5017 (.I0(STAGE4_EN), .I1(n221), .O(n30807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5017.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5018 (.I0(\ARG2[11] ), .I1(\ARG1[11] ), .I2(\ARG2[12] ), 
            .I3(\ARG1[12] ), .O(n3446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5018.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5019 (.I0(\ARG1[12] ), .I1(\ARG2[12] ), .O(n3447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5019.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5020 (.I0(\ARG2[6] ), .I1(\ARG1[6] ), .I2(\ARG2[7] ), 
            .I3(\ARG1[7] ), .O(n3448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5020.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5021 (.I0(\ARG1[7] ), .I1(\ARG2[7] ), .I2(\ARG1[8] ), 
            .I3(\ARG2[8] ), .O(n3449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5021.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5022 (.I0(\ARG2[10] ), .I1(\ARG1[10] ), .O(n3450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5022.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5023 (.I0(\ARG2[8] ), .I1(\ARG1[8] ), .I2(\ARG2[9] ), 
            .I3(\ARG1[9] ), .O(n3451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5023.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5024 (.I0(n3449), .I1(n3448), .I2(n3450), .I3(n3451), 
            .O(n3452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__5024.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__5025 (.I0(\ARG2[10] ), .I1(\ARG1[10] ), .I2(\ARG1[9] ), 
            .I3(\ARG2[9] ), .O(n3453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__5025.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__5026 (.I0(\ARG2[11] ), .I1(\ARG1[11] ), .I2(n3447), 
            .I3(n3453), .O(n3454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__5026.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__5027 (.I0(n3452), .I1(n3454), .I2(n3446), .I3(n3447), 
            .O(n3455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__5027.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__5028 (.I0(\ARG1[1] ), .I1(\ARG1[0] ), .I2(\ARG2[0] ), 
            .I3(\ARG2[1] ), .O(n3456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5028.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5029 (.I0(\ARG1[0] ), .I1(\ARG2[0] ), .I2(\ARG1[1] ), 
            .O(n3457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__5029.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__5030 (.I0(\ARG2[4] ), .I1(\ARG1[4] ), .I2(\ARG2[5] ), 
            .I3(\ARG1[5] ), .O(n3458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5030.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5031 (.I0(\ARG2[3] ), .I1(\ARG1[3] ), .I2(\ARG2[2] ), 
            .I3(\ARG1[2] ), .O(n3459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5031.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5032 (.I0(n3456), .I1(n3457), .I2(n3458), .I3(n3459), 
            .O(n3460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5032.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5033 (.I0(\ARG1[2] ), .I1(\ARG2[2] ), .O(n3461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5033.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5034 (.I0(n3461), .I1(\ARG1[3] ), .I2(\ARG2[3] ), .I3(n3458), 
            .O(n3462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__5034.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__5035 (.I0(\ARG1[6] ), .I1(\ARG2[6] ), .O(n3463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5035.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5036 (.I0(\ARG2[5] ), .I1(\ARG1[5] ), .I2(\ARG1[4] ), 
            .I3(\ARG2[4] ), .O(n3464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__5036.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__5037 (.I0(n3463), .I1(n3464), .I2(n3449), .O(n3465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5037.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5038 (.I0(n3460), .I1(n3462), .I2(n3465), .I3(n3454), 
            .O(n3466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5038.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5039 (.I0(\ARG2[16] ), .I1(\ARG1[16] ), .I2(\ARG1[15] ), 
            .I3(\ARG2[15] ), .O(n3467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__5039.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__5040 (.I0(\ARG1[17] ), .I1(\ARG2[17] ), .I2(\ARG1[18] ), 
            .I3(\ARG2[18] ), .O(n3468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5040.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5041 (.I0(n3467), .I1(n3468), .O(n3469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5041.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5042 (.I0(\ARG1[14] ), .I1(\ARG2[14] ), .O(n3470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5042.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5043 (.I0(n3470), .I1(\ARG1[13] ), .O(n3471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5043.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5044 (.I0(n3466), .I1(n3455), .I2(n3469), .I3(n3471), 
            .O(n3472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__5044.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__5045 (.I0(\ARG2[14] ), .I1(\ARG1[14] ), .I2(\ARG2[15] ), 
            .I3(\ARG1[15] ), .O(n3473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5045.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5046 (.I0(\ARG2[16] ), .I1(\ARG1[16] ), .I2(n3473), 
            .O(n3474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__5046.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__5047 (.I0(\ARG1[13] ), .I1(n3446), .O(n3475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5047.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5048 (.I0(n3452), .I1(n3474), .I2(n3475), .O(n3476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__5048.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__5049 (.I0(n3460), .I1(n3462), .I2(n3465), .O(n3477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5049.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5050 (.I0(\ARG2[12] ), .I1(\ARG1[12] ), .I2(\ARG1[11] ), 
            .I3(\ARG2[11] ), .O(n3478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__5050.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__5051 (.I0(n3478), .I1(\ARG1[13] ), .I2(\ARG2[13] ), 
            .I3(n3470), .O(n3479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__5051.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__5052 (.I0(n3453), .I1(n3475), .I2(n3479), .I3(n3474), 
            .O(n3480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__5052.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__5053 (.I0(n3477), .I1(n3476), .I2(n3480), .I3(n3469), 
            .O(n3481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__5053.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__5054 (.I0(\ARG2[22] ), .I1(\ARG1[22] ), .O(n3482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5054.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5055 (.I0(\ARG2[21] ), .I1(\ARG2[20] ), .I2(\ARG1[21] ), 
            .I3(\ARG1[20] ), .O(n3483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__5055.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__5056 (.I0(\ARG1[23] ), .I1(\ARG2[23] ), .I2(\ARG1[22] ), 
            .I3(\ARG2[22] ), .O(n3484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5056.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5057 (.I0(\ARG2[23] ), .I1(\ARG1[23] ), .O(n3485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5057.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5058 (.I0(n3482), .I1(n3483), .I2(n3484), .I3(n3485), 
            .O(n3486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5058.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5059 (.I0(\ARG2[25] ), .I1(\ARG1[25] ), .I2(\ARG2[24] ), 
            .I3(\ARG1[24] ), .O(n3487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5059.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5060 (.I0(\ARG2[26] ), .I1(\ARG1[26] ), .I2(n3487), 
            .O(n3488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__5060.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__5061 (.I0(\ARG2[18] ), .I1(\ARG2[17] ), .I2(\ARG1[18] ), 
            .I3(\ARG1[17] ), .O(n3489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__5061.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__5062 (.I0(\ARG2[19] ), .I1(\ARG1[19] ), .I2(n3489), 
            .O(n3490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__5062.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__5063 (.I0(n3486), .I1(n3488), .I2(n3490), .O(n3491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__5063.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__5064 (.I0(\ARG2[29] ), .I1(\ARG1[29] ), .I2(\ARG2[28] ), 
            .I3(\ARG1[28] ), .O(n3492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5064.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5065 (.I0(\ARG1[27] ), .I1(\ARG2[27] ), .I2(n3492), 
            .O(n3493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5065.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5066 (.I0(n3491), .I1(n3493), .O(n3494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5066.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5067 (.I0(\ARG1[19] ), .I1(\ARG2[19] ), .I2(\ARG1[20] ), 
            .I3(\ARG2[20] ), .O(n3495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5067.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5068 (.I0(\ARG2[21] ), .I1(\ARG1[21] ), .I2(n3484), 
            .I3(n3495), .O(n3496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__5068.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__5069 (.I0(\ARG2[25] ), .I1(\ARG1[25] ), .I2(\ARG1[24] ), 
            .I3(\ARG2[24] ), .O(n3497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__5069.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__5070 (.I0(n3497), .I1(\ARG1[26] ), .I2(\ARG2[26] ), 
            .O(n3498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__5070.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__5071 (.I0(n3496), .I1(n3486), .I2(n3488), .I3(n3498), 
            .O(n3499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__5071.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__5072 (.I0(\ARG1[28] ), .I1(\ARG2[28] ), .I2(\ARG1[27] ), 
            .I3(\ARG2[27] ), .O(n3500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5072.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5073 (.I0(n3500), .I1(n3492), .I2(\ARG1[29] ), .I3(\ARG2[29] ), 
            .O(n3501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__5073.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__5074 (.I0(n3499), .I1(n3493), .I2(n3501), .O(n3502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__5074.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__5075 (.I0(n3481), .I1(n3472), .I2(n3494), .I3(n3502), 
            .O(n2741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5075.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5076 (.I0(\ARG2[31] ), .I1(\ARG1[31] ), .O(n3503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__5076.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__5077 (.I0(\ARG2[30] ), .I1(\ARG1[30] ), .I2(n3503), 
            .I3(\OPERATION[3] ), .O(n3504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__5077.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__5078 (.I0(\ARG1[7] ), .I1(\ARG1[5] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5078.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5079 (.I0(\ARG1[6] ), .I1(\ARG1[4] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5079.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5080 (.I0(n3506), .I1(n3505), .I2(\SHIFT_STEPS[0] ), 
            .O(n3507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5080.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5081 (.I0(\SHIFT_STEPS[1] ), .I1(\ARG1[1] ), .O(n3508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5081.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5082 (.I0(\SHIFT_STEPS[1] ), .I1(\ARG1[3] ), .O(n3509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5082.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5083 (.I0(\ARG1[0] ), .I1(\ARG1[2] ), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[1] ), .O(n3510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5083.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5084 (.I0(n3509), .I1(n3508), .I2(\SHIFT_STEPS[0] ), 
            .I3(n3510), .O(n3511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5084.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5085 (.I0(n3511), .I1(n3507), .I2(\SHIFT_STEPS[2] ), 
            .O(n3512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5085.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5086 (.I0(\ARG1[15] ), .I1(\ARG1[13] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5086.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5087 (.I0(\ARG1[14] ), .I1(\ARG1[12] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5087.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5088 (.I0(n3514), .I1(n3513), .I2(\SHIFT_STEPS[0] ), 
            .O(n3515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5088.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5089 (.I0(\ARG1[11] ), .I1(\ARG1[9] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5089.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5090 (.I0(\ARG1[10] ), .I1(\ARG1[8] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5090.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5091 (.I0(n3517), .I1(n3516), .I2(\SHIFT_STEPS[0] ), 
            .O(n3518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5091.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5092 (.I0(n3518), .I1(n3515), .I2(\SHIFT_STEPS[2] ), 
            .O(n3519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__5092.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__5093 (.I0(n3519), .I1(n3512), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n3520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__5093.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__5094 (.I0(\ARG1[31] ), .I1(\ARG1[29] ), .I2(\SHIFT_STEPS[1] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n3521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__5094.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__5095 (.I0(\ARG1[30] ), .I1(\ARG1[28] ), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[1] ), .O(n3522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5095.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5096 (.I0(n3521), .I1(n3522), .O(n3523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5096.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5097 (.I0(\ARG1[27] ), .I1(\ARG1[25] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5097.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5098 (.I0(\ARG1[26] ), .I1(\ARG1[24] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5098.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5099 (.I0(n3525), .I1(n3524), .I2(\SHIFT_STEPS[0] ), 
            .O(n3526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5099.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5100 (.I0(n3526), .I1(n3523), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n3527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__5100.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__5101 (.I0(\ARG1[23] ), .I1(\ARG1[21] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5101.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5102 (.I0(\ARG1[22] ), .I1(\ARG1[20] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5102.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5103 (.I0(n3529), .I1(n3528), .I2(\SHIFT_STEPS[0] ), 
            .O(n3530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5103.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5104 (.I0(\ARG1[19] ), .I1(\ARG1[17] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5104.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5105 (.I0(\ARG1[18] ), .I1(\ARG1[16] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n3532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5105.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5106 (.I0(n3532), .I1(n3531), .I2(\SHIFT_STEPS[0] ), 
            .O(n3533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5106.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5107 (.I0(n3533), .I1(n3530), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n3534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5107.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5108 (.I0(n3534), .I1(n3527), .I2(\SHIFT_STEPS[4] ), 
            .O(n3535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__5108.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__5109 (.I0(\OPERATION[0] ), .I1(\OPERATION[1] ), .O(n3536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5109.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5110 (.I0(\OPERATION[3] ), .I1(\OPERATION[2] ), .O(n3537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5110.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5111 (.I0(\OPERATION[0] ), .I1(\ARG1[0] ), .I2(\OPERATION[1] ), 
            .I3(\ARG2[0] ), .O(n3538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__5111.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__5112 (.I0(n3537), .I1(n3538), .O(n3539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5112.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5113 (.I0(n3535), .I1(n3520), .I2(n3536), .I3(n3539), 
            .O(n3540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__5113.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__5114 (.I0(\SHIFT_STEPS[0] ), .I1(\SHIFT_STEPS[1] ), .I2(\ARG1[0] ), 
            .O(n3541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5114.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5115 (.I0(\SHIFT_STEPS[2] ), .I1(\SHIFT_STEPS[3] ), .O(n3542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5115.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5116 (.I0(\SHIFT_STEPS[4] ), .I1(n3542), .I2(n3445), 
            .O(n3543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5116.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5117 (.I0(n8), .I1(n39), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n3544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5117.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5118 (.I0(\OPERATION[2] ), .I1(\OPERATION[3] ), .O(n3545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5118.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5119 (.I0(n3543), .I1(n3541), .I2(n3544), .I3(n3545), 
            .O(n3546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__5119.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__5120 (.I0(\OPERATION[0] ), .I1(\OPERATION[1] ), .O(n3547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5120.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5121 (.I0(\OPERATION[3] ), .I1(\OPERATION[0] ), .I2(\ARG2[31] ), 
            .I3(\ARG1[31] ), .O(n3548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha82a */ ;
    defparam LUT__5121.LUTMASK = 16'ha82a;
    EFX_LUT4 LUT__5122 (.I0(\ARG1[30] ), .I1(\ARG2[30] ), .I2(n3503), 
            .I3(n3548), .O(n3549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__5122.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__5123 (.I0(n3546), .I1(n3547), .I2(n3549), .O(n3550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__5123.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__5124 (.I0(n3535), .I1(n3520), .I2(n3546), .I3(n3550), 
            .O(n3551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5124.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5125 (.I0(\RES[0]_2~FF_brt_192_q ), .I1(\RES[0]_2~FF_brt_193_q ), 
            .I2(\RES[0]_2~FF_brt_194_q ), .I3(\RES[0]_2~FF_brt_195_q ), 
            .O(n1615_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5125.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5126 (.I0(\OPERATION[1] ), .I1(\OPERATION[2] ), .O(n3552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5126.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5127 (.I0(n3552), .I1(\OPERATION[3] ), .I2(n30678), 
            .O(ceg_net408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__5127.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__5128 (.I0(STAGE2_EN), .I1(n51814), .O(\INSTRUCTION[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5128.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5129 (.I0(STAGE2_EN), .I1(n51810), .O(\INSTRUCTION[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5129.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5130 (.I0(STAGE2_EN), .I1(n51806), .O(\INSTRUCTION[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5130.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5131 (.I0(STAGE2_EN), .I1(n51750), .O(\INSTRUCTION[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5131.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5132 (.I0(STAGE2_EN), .I1(n51746), .O(\INSTRUCTION[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5132.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5133 (.I0(STAGE2_EN), .I1(n51742), .O(\INSTRUCTION[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5133.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5134 (.I0(STAGE2_EN), .I1(n51738), .O(\INSTRUCTION[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5134.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5135 (.I0(STAGE2_EN), .I1(n51734), .O(\INSTRUCTION[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5135.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5136 (.I0(n3547), .I1(\OPERATION[3] ), .O(n34248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5136.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5137 (.I0(n3145), .I1(n2953), .I2(n3203), .O(n540_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__5137.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__5138 (.I0(n3087), .I1(n2959), .I2(n3203), .O(n539_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__5138.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__5139 (.I0(n3058), .I1(n2967), .I2(n3203), .O(n538_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5139.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5140 (.I0(n3203), .I1(n2966), .O(n537_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5140.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5141 (.I0(n51802), .I1(n51794), .O(n3553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5141.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5142 (.I0(n51730), .I1(n51794), .I2(n51798), .I3(n51802), 
            .O(n3554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__5142.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__5143 (.I0(n3554), .I1(n3553), .I2(n2982), .I3(n3202), 
            .O(n530_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5143.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5144 (.I0(n3202), .I1(n3554), .I2(n2982), .I3(n51794), 
            .O(n529_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5144.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5145 (.I0(n51794), .I1(n51798), .I2(n2982), .I3(n3202), 
            .O(n528_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5145.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5146 (.I0(n51798), .I1(n51830), .I2(n51802), .I3(n51794), 
            .O(n3555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3001 */ ;
    defparam LUT__5146.LUTMASK = 16'h3001;
    EFX_LUT4 LUT__5147 (.I0(\DATA_FORMAT[1] ), .I1(n51830), .I2(n51798), 
            .I3(n51802), .O(n3556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__5147.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__5148 (.I0(n3555), .I1(n3556), .I2(STAGE2_EN), .O(n33468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__5148.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__5149 (.I0(n51798), .I1(n51802), .I2(\DATA_FORMAT[2] ), 
            .I3(n3208), .O(n3557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5149.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5150 (.I0(n3557), .I1(n3553), .I2(n51830), .I3(STAGE2_EN), 
            .O(n33460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__5150.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__5151 (.I0(n3208), .I1(STAGE2_EN), .I2(n51802), .I3(n51798), 
            .O(n3558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__5151.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__5152 (.I0(n3558), .I1(n3211), .O(ceg_net47657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__5152.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__5153 (.I0(STAGE2_EN), .I1(n51818), .O(\INSTRUCTION[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5153.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5154 (.I0(n34248), .I1(n30678), .O(n50605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5154.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5155 (.I0(\DATA_FORMAT_2[2] ), .I1(\DATA_FORMAT_2[0] ), 
            .I2(\DATA_FORMAT_2[1] ), .I3(n50605), .O(ceg_net35302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4300 */ ;
    defparam LUT__5155.LUTMASK = 16'h4300;
    EFX_LUT4 LUT__5156 (.I0(\XI[18][14] ), .I1(\XI[19][14] ), .I2(n51770), 
            .O(n3559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5156.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5157 (.I0(\XI[16][14] ), .I1(\XI[17][14] ), .I2(n51770), 
            .O(n3560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5157.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5158 (.I0(n3559), .I1(n3560), .I2(n2959), .I3(n2953), 
            .O(n3561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5158.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5159 (.I0(\XI[21][14] ), .I1(\XI[20][14] ), .I2(n2953), 
            .I3(n2954), .O(n3562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5159.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5160 (.I0(\XI[23][14] ), .I1(\XI[22][14] ), .I2(n51770), 
            .O(n3563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5160.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5161 (.I0(n3563), .I1(n3561), .I2(n3562), .I3(n2959), 
            .O(n3564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5161.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5162 (.I0(\XI[25][14] ), .I1(\XI[24][14] ), .I2(n2954), 
            .O(n3565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5162.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5163 (.I0(\XI[27][14] ), .I1(\XI[26][14] ), .I2(n2954), 
            .O(n3566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5163.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5164 (.I0(n3566), .I1(n3565), .I2(n2959), .I3(n2953), 
            .O(n3567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5164.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5165 (.I0(\XI[31][14] ), .I1(\XI[30][14] ), .I2(n2954), 
            .O(n3568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5165.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5166 (.I0(\XI[29][14] ), .I1(\XI[28][14] ), .I2(n2954), 
            .O(n3569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5166.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5167 (.I0(n3569), .I1(n3568), .I2(n2953), .I3(n2959), 
            .O(n3570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5167.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5168 (.I0(n3567), .I1(n3570), .I2(n3564), .I3(n2967), 
            .O(n3571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5168.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5169 (.I0(\XI[15][14] ), .I1(\XI[14][14] ), .I2(n2954), 
            .I3(n2953), .O(n3572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5169.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5170 (.I0(\XI[13][14] ), .I1(\XI[12][14] ), .I2(n2953), 
            .I3(n2954), .O(n3573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5170.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5171 (.I0(n3572), .I1(n3573), .I2(n2959), .O(n3574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5171.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5172 (.I0(\XI[9][14] ), .I1(\XI[8][14] ), .I2(n2954), 
            .O(n3575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5172.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5173 (.I0(\XI[11][14] ), .I1(\XI[10][14] ), .I2(n2954), 
            .O(n3576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5173.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5174 (.I0(n3576), .I1(n3575), .I2(n2959), .I3(n2953), 
            .O(n3577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5174.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5175 (.I0(\XI[5][14] ), .I1(\XI[4][14] ), .I2(n2953), 
            .I3(n2954), .O(n3578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5175.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5176 (.I0(\XI[7][14] ), .I1(\XI[6][14] ), .I2(n2954), 
            .I3(n2953), .O(n3579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5176.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5180 (.I0(n3579), .I1(n3578), .I2(n3582), .I3(n2959), 
            .O(n3583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5180.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5181 (.I0(n3577), .I1(n3574), .I2(n3583), .I3(n2967), 
            .O(n3584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5181.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5182 (.I0(n3584), .I1(n3571), .I2(n3029), .I3(n2966), 
            .O(n3585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5182.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5183 (.I0(\PC[14] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5183.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5184 (.I0(n3584), .I1(n3571), .I2(n2991), .I3(n2966), 
            .O(n3587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5184.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5185 (.I0(n2983), .I1(\PC[14] ), .I2(n3383), .O(n3588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5185.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5186 (.I0(n3587), .I1(n3588), .I2(n3585), .I3(n3586), 
            .O(n512_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5186.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5187 (.I0(\XI[18][15] ), .I1(\XI[19][15] ), .I2(n51770), 
            .O(n3589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5187.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5188 (.I0(\XI[16][15] ), .I1(\XI[17][15] ), .I2(n51770), 
            .O(n3590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5188.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5189 (.I0(n3589), .I1(n3590), .I2(n2959), .I3(n2953), 
            .O(n3591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5189.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5190 (.I0(\XI[21][15] ), .I1(\XI[20][15] ), .I2(n2953), 
            .I3(n2954), .O(n3592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5190.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5191 (.I0(\XI[23][15] ), .I1(\XI[22][15] ), .I2(n51770), 
            .O(n3593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5191.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5192 (.I0(n3593), .I1(n3591), .I2(n3592), .I3(n2959), 
            .O(n3594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5192.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5193 (.I0(\XI[25][15] ), .I1(\XI[24][15] ), .I2(n2954), 
            .O(n3595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5193.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5194 (.I0(\XI[27][15] ), .I1(\XI[26][15] ), .I2(n2954), 
            .O(n3596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5194.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5195 (.I0(n3596), .I1(n3595), .I2(n2959), .I3(n2953), 
            .O(n3597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5195.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5196 (.I0(\XI[31][15] ), .I1(\XI[30][15] ), .I2(n2954), 
            .O(n3598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5196.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5197 (.I0(\XI[29][15] ), .I1(\XI[28][15] ), .I2(n2954), 
            .O(n3599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5197.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5198 (.I0(n3599), .I1(n3598), .I2(n2953), .I3(n2959), 
            .O(n3600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5198.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5199 (.I0(n3597), .I1(n3600), .I2(n3594), .I3(n2967), 
            .O(n3601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5199.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5200 (.I0(\XI[15][15] ), .I1(\XI[14][15] ), .I2(n2954), 
            .I3(n2953), .O(n3602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5200.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5201 (.I0(\XI[13][15] ), .I1(\XI[12][15] ), .I2(n2953), 
            .I3(n2954), .O(n3603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5201.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5202 (.I0(n3602), .I1(n3603), .I2(n2959), .O(n3604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5202.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5203 (.I0(\XI[9][15] ), .I1(\XI[8][15] ), .I2(n2954), 
            .O(n3605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5203.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5204 (.I0(\XI[11][15] ), .I1(\XI[10][15] ), .I2(n2954), 
            .O(n3606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5204.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5205 (.I0(n3606), .I1(n3605), .I2(n2959), .I3(n2953), 
            .O(n3607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5205.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5206 (.I0(\XI[5][15] ), .I1(\XI[4][15] ), .I2(n2953), 
            .I3(n2954), .O(n3608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5206.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5207 (.I0(\XI[7][15] ), .I1(\XI[6][15] ), .I2(n2954), 
            .I3(n2953), .O(n3609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5207.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5211 (.I0(n3609), .I1(n3608), .I2(n3612), .I3(n2959), 
            .O(n3613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5211.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5212 (.I0(n3607), .I1(n3604), .I2(n3613), .I3(n2967), 
            .O(n3614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5212.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5213 (.I0(n3614), .I1(n3601), .I2(n3029), .I3(n2966), 
            .O(n3615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5213.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5214 (.I0(\PC[15] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5214.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5215 (.I0(n3614), .I1(n3601), .I2(n2991), .I3(n2966), 
            .O(n3617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5215.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5216 (.I0(n2983), .I1(\PC[15] ), .I2(n3383), .O(n3618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5216.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5217 (.I0(n3617), .I1(n3618), .I2(n3615), .I3(n3616), 
            .O(n511_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5217.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5218 (.I0(\XI[18][16] ), .I1(\XI[19][16] ), .I2(n51770), 
            .O(n3619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5218.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5219 (.I0(\XI[16][16] ), .I1(\XI[17][16] ), .I2(n51770), 
            .O(n3620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5219.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5220 (.I0(n3619), .I1(n3620), .I2(n2959), .I3(n2953), 
            .O(n3621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5220.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5221 (.I0(\XI[21][16] ), .I1(\XI[20][16] ), .I2(n2953), 
            .I3(n2954), .O(n3622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5221.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5222 (.I0(\XI[23][16] ), .I1(\XI[22][16] ), .I2(n51770), 
            .O(n3623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5222.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5223 (.I0(n3623), .I1(n3621), .I2(n3622), .I3(n2959), 
            .O(n3624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5223.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5224 (.I0(\XI[25][16] ), .I1(\XI[24][16] ), .I2(n2954), 
            .O(n3625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5224.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5225 (.I0(\XI[27][16] ), .I1(\XI[26][16] ), .I2(n2954), 
            .O(n3626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5225.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5226 (.I0(n3626), .I1(n3625), .I2(n2959), .I3(n2953), 
            .O(n3627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5226.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5227 (.I0(\XI[31][16] ), .I1(\XI[30][16] ), .I2(n2954), 
            .O(n3628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5227.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5228 (.I0(\XI[29][16] ), .I1(\XI[28][16] ), .I2(n2954), 
            .O(n3629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5228.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5229 (.I0(n3629), .I1(n3628), .I2(n2953), .I3(n2959), 
            .O(n3630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5229.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5230 (.I0(n3627), .I1(n3630), .I2(n3624), .I3(n2967), 
            .O(n3631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5230.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5231 (.I0(\XI[15][16] ), .I1(\XI[14][16] ), .I2(n2954), 
            .I3(n2953), .O(n3632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5231.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5232 (.I0(\XI[13][16] ), .I1(\XI[12][16] ), .I2(n2953), 
            .I3(n2954), .O(n3633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5232.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5233 (.I0(n3632), .I1(n3633), .I2(n2959), .O(n3634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5233.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5234 (.I0(\XI[9][16] ), .I1(\XI[8][16] ), .I2(n2954), 
            .O(n3635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5234.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5235 (.I0(\XI[11][16] ), .I1(\XI[10][16] ), .I2(n2954), 
            .O(n3636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5235.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5236 (.I0(n3636), .I1(n3635), .I2(n2959), .I3(n2953), 
            .O(n3637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5236.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5237 (.I0(\XI[5][16] ), .I1(\XI[4][16] ), .I2(n2953), 
            .I3(n2954), .O(n3638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5237.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5238 (.I0(\XI[7][16] ), .I1(\XI[6][16] ), .I2(n2954), 
            .I3(n2953), .O(n3639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5238.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5242 (.I0(n3639), .I1(n3638), .I2(n3642), .I3(n2959), 
            .O(n3643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5242.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5243 (.I0(n3637), .I1(n3634), .I2(n3643), .I3(n2967), 
            .O(n3644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5243.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5244 (.I0(n3644), .I1(n3631), .I2(n3029), .I3(n2966), 
            .O(n3645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5244.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5245 (.I0(\PC[16] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5245.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5246 (.I0(n3644), .I1(n3631), .I2(n2991), .I3(n2966), 
            .O(n3647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5246.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5247 (.I0(n2983), .I1(\PC[16] ), .I2(n3383), .O(n3648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5247.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5248 (.I0(n3647), .I1(n3648), .I2(n3645), .I3(n3646), 
            .O(n510_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5248.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5249 (.I0(\XI[18][17] ), .I1(\XI[19][17] ), .I2(n51770), 
            .O(n3649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5249.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5250 (.I0(\XI[16][17] ), .I1(\XI[17][17] ), .I2(n51770), 
            .O(n3650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5250.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5251 (.I0(n3649), .I1(n3650), .I2(n2959), .I3(n2953), 
            .O(n3651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5251.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5252 (.I0(\XI[21][17] ), .I1(\XI[20][17] ), .I2(n2953), 
            .I3(n2954), .O(n3652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5252.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5253 (.I0(\XI[23][17] ), .I1(\XI[22][17] ), .I2(n51770), 
            .O(n3653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5253.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5254 (.I0(n3653), .I1(n3651), .I2(n3652), .I3(n2959), 
            .O(n3654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5254.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5255 (.I0(\XI[25][17] ), .I1(\XI[24][17] ), .I2(n2954), 
            .O(n3655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5255.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5256 (.I0(\XI[27][17] ), .I1(\XI[26][17] ), .I2(n2954), 
            .O(n3656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5256.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5257 (.I0(n3656), .I1(n3655), .I2(n2959), .I3(n2953), 
            .O(n3657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5257.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5258 (.I0(\XI[31][17] ), .I1(\XI[30][17] ), .I2(n2954), 
            .O(n3658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5258.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5259 (.I0(\XI[29][17] ), .I1(\XI[28][17] ), .I2(n2954), 
            .O(n3659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5259.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5260 (.I0(n3659), .I1(n3658), .I2(n2953), .I3(n2959), 
            .O(n3660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5260.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5261 (.I0(n3657), .I1(n3660), .I2(n3654), .I3(n2967), 
            .O(n3661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5261.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5262 (.I0(\XI[15][17] ), .I1(\XI[14][17] ), .I2(n2954), 
            .I3(n2953), .O(n3662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5262.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5263 (.I0(\XI[13][17] ), .I1(\XI[12][17] ), .I2(n2953), 
            .I3(n2954), .O(n3663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5263.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5264 (.I0(n3662), .I1(n3663), .I2(n2959), .O(n3664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5264.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5265 (.I0(\XI[9][17] ), .I1(\XI[8][17] ), .I2(n2954), 
            .O(n3665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5265.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5266 (.I0(\XI[11][17] ), .I1(\XI[10][17] ), .I2(n2954), 
            .O(n3666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5266.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5267 (.I0(n3666), .I1(n3665), .I2(n2959), .I3(n2953), 
            .O(n3667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5267.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5268 (.I0(\XI[5][17] ), .I1(\XI[4][17] ), .I2(n2953), 
            .I3(n2954), .O(n3668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5268.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5269 (.I0(\XI[7][17] ), .I1(\XI[6][17] ), .I2(n2954), 
            .I3(n2953), .O(n3669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5269.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5273 (.I0(n3669), .I1(n3668), .I2(n3672), .I3(n2959), 
            .O(n3673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5273.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5274 (.I0(n3667), .I1(n3664), .I2(n3673), .I3(n2967), 
            .O(n3674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5274.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5275 (.I0(n3674), .I1(n3661), .I2(n3029), .I3(n2966), 
            .O(n3675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5275.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5276 (.I0(\PC[17] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5276.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5277 (.I0(n3674), .I1(n3661), .I2(n2991), .I3(n2966), 
            .O(n3677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5277.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5278 (.I0(n2983), .I1(\PC[17] ), .I2(n3383), .O(n3678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5278.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5279 (.I0(n3677), .I1(n3678), .I2(n3675), .I3(n3676), 
            .O(n509_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5279.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5280 (.I0(\XI[18][18] ), .I1(\XI[19][18] ), .I2(n51770), 
            .O(n3679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5280.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5281 (.I0(\XI[16][18] ), .I1(\XI[17][18] ), .I2(n51770), 
            .O(n3680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5281.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5282 (.I0(n3679), .I1(n3680), .I2(n2959), .I3(n2953), 
            .O(n3681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5282.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5283 (.I0(\XI[21][18] ), .I1(\XI[20][18] ), .I2(n2953), 
            .I3(n2954), .O(n3682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5283.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5284 (.I0(\XI[23][18] ), .I1(\XI[22][18] ), .I2(n51770), 
            .O(n3683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5284.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5285 (.I0(n3683), .I1(n3681), .I2(n3682), .I3(n2959), 
            .O(n3684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5285.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5286 (.I0(\XI[25][18] ), .I1(\XI[24][18] ), .I2(n2954), 
            .O(n3685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5286.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5287 (.I0(\XI[27][18] ), .I1(\XI[26][18] ), .I2(n2954), 
            .O(n3686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5287.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5288 (.I0(n3686), .I1(n3685), .I2(n2959), .I3(n2953), 
            .O(n3687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5288.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5289 (.I0(\XI[31][18] ), .I1(\XI[30][18] ), .I2(n2954), 
            .O(n3688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5289.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5290 (.I0(\XI[29][18] ), .I1(\XI[28][18] ), .I2(n2954), 
            .O(n3689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5290.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5291 (.I0(n3689), .I1(n3688), .I2(n2953), .I3(n2959), 
            .O(n3690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5291.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5292 (.I0(n3687), .I1(n3690), .I2(n3684), .I3(n2967), 
            .O(n3691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5292.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5293 (.I0(\XI[15][18] ), .I1(\XI[14][18] ), .I2(n2954), 
            .I3(n2953), .O(n3692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5293.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5294 (.I0(\XI[13][18] ), .I1(\XI[12][18] ), .I2(n2953), 
            .I3(n2954), .O(n3693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5294.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5295 (.I0(n3692), .I1(n3693), .I2(n2959), .O(n3694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5295.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5296 (.I0(\XI[9][18] ), .I1(\XI[8][18] ), .I2(n2954), 
            .O(n3695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5296.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5297 (.I0(\XI[11][18] ), .I1(\XI[10][18] ), .I2(n2954), 
            .O(n3696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5297.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5298 (.I0(n3696), .I1(n3695), .I2(n2959), .I3(n2953), 
            .O(n3697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5298.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5299 (.I0(\XI[5][18] ), .I1(\XI[4][18] ), .I2(n2953), 
            .I3(n2954), .O(n3698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5299.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5300 (.I0(\XI[7][18] ), .I1(\XI[6][18] ), .I2(n2954), 
            .I3(n2953), .O(n3699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5300.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5304 (.I0(n3699), .I1(n3698), .I2(n3702), .I3(n2959), 
            .O(n3703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5304.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5305 (.I0(n3697), .I1(n3694), .I2(n3703), .I3(n2967), 
            .O(n3704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5305.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5306 (.I0(n3704), .I1(n3691), .I2(n3029), .I3(n2966), 
            .O(n3705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5306.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5307 (.I0(\PC[18] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5307.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5308 (.I0(n3704), .I1(n3691), .I2(n2991), .I3(n2966), 
            .O(n3707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5308.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5309 (.I0(n2983), .I1(\PC[18] ), .I2(n3383), .O(n3708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5309.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5310 (.I0(n3707), .I1(n3708), .I2(n3705), .I3(n3706), 
            .O(n508_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5310.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5311 (.I0(\XI[18][19] ), .I1(\XI[19][19] ), .I2(n51770), 
            .O(n3709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5311.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5312 (.I0(\XI[16][19] ), .I1(\XI[17][19] ), .I2(n51770), 
            .O(n3710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5312.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5313 (.I0(n3709), .I1(n3710), .I2(n2959), .I3(n2953), 
            .O(n3711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5313.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5314 (.I0(\XI[21][19] ), .I1(\XI[20][19] ), .I2(n2953), 
            .I3(n2954), .O(n3712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5314.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5315 (.I0(\XI[23][19] ), .I1(\XI[22][19] ), .I2(n51770), 
            .O(n3713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5315.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5316 (.I0(n3713), .I1(n3711), .I2(n3712), .I3(n2959), 
            .O(n3714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5316.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5317 (.I0(\XI[25][19] ), .I1(\XI[24][19] ), .I2(n2954), 
            .O(n3715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5317.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5318 (.I0(\XI[27][19] ), .I1(\XI[26][19] ), .I2(n2954), 
            .O(n3716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5318.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5319 (.I0(n3716), .I1(n3715), .I2(n2959), .I3(n2953), 
            .O(n3717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5319.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5320 (.I0(\XI[31][19] ), .I1(\XI[30][19] ), .I2(n2954), 
            .O(n3718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5320.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5321 (.I0(\XI[29][19] ), .I1(\XI[28][19] ), .I2(n2954), 
            .O(n3719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5321.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5322 (.I0(n3719), .I1(n3718), .I2(n2953), .I3(n2959), 
            .O(n3720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5322.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5323 (.I0(n3717), .I1(n3720), .I2(n3714), .I3(n2967), 
            .O(n3721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5323.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5324 (.I0(\XI[15][19] ), .I1(\XI[14][19] ), .I2(n2954), 
            .I3(n2953), .O(n3722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5324.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5325 (.I0(\XI[13][19] ), .I1(\XI[12][19] ), .I2(n2953), 
            .I3(n2954), .O(n3723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5325.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5326 (.I0(n3722), .I1(n3723), .I2(n2959), .O(n3724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5326.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5327 (.I0(\XI[9][19] ), .I1(\XI[8][19] ), .I2(n2954), 
            .O(n3725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5327.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5328 (.I0(\XI[11][19] ), .I1(\XI[10][19] ), .I2(n2954), 
            .O(n3726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5328.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5329 (.I0(n3726), .I1(n3725), .I2(n2959), .I3(n2953), 
            .O(n3727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5329.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5330 (.I0(\XI[5][19] ), .I1(\XI[4][19] ), .I2(n2953), 
            .I3(n2954), .O(n3728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5330.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5331 (.I0(\XI[7][19] ), .I1(\XI[6][19] ), .I2(n2954), 
            .I3(n2953), .O(n3729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5331.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5335 (.I0(n3729), .I1(n3728), .I2(n3732), .I3(n2959), 
            .O(n3733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5335.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5336 (.I0(n3727), .I1(n3724), .I2(n3733), .I3(n2967), 
            .O(n3734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5336.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5337 (.I0(n3734), .I1(n3721), .I2(n3029), .I3(n2966), 
            .O(n3735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5337.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5338 (.I0(\PC[19] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5338.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5339 (.I0(n3734), .I1(n3721), .I2(n2991), .I3(n2966), 
            .O(n3737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5339.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5340 (.I0(n2983), .I1(\PC[19] ), .I2(n3383), .O(n3738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5340.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5341 (.I0(n3737), .I1(n3738), .I2(n3735), .I3(n3736), 
            .O(n507_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5341.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5342 (.I0(\XI[18][25] ), .I1(\XI[19][25] ), .I2(n51770), 
            .O(n3739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5342.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5343 (.I0(\XI[16][25] ), .I1(\XI[17][25] ), .I2(n51770), 
            .O(n3740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5343.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5344 (.I0(n3739), .I1(n3740), .I2(n2959), .I3(n2953), 
            .O(n3741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5344.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5345 (.I0(\XI[21][25] ), .I1(\XI[20][25] ), .I2(n2953), 
            .I3(n2954), .O(n3742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5345.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5346 (.I0(\XI[23][25] ), .I1(\XI[22][25] ), .I2(n51770), 
            .O(n3743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5346.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5347 (.I0(n3743), .I1(n3741), .I2(n3742), .I3(n2959), 
            .O(n3744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5347.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5348 (.I0(\XI[25][25] ), .I1(\XI[24][25] ), .I2(n2954), 
            .O(n3745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5348.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5349 (.I0(\XI[27][25] ), .I1(\XI[26][25] ), .I2(n2954), 
            .O(n3746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5349.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5350 (.I0(n3746), .I1(n3745), .I2(n2959), .I3(n2953), 
            .O(n3747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5350.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5351 (.I0(\XI[31][25] ), .I1(\XI[30][25] ), .I2(n2954), 
            .O(n3748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5351.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5352 (.I0(\XI[29][25] ), .I1(\XI[28][25] ), .I2(n2954), 
            .O(n3749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5352.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5353 (.I0(n3749), .I1(n3748), .I2(n2953), .I3(n2959), 
            .O(n3750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5353.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5354 (.I0(n3747), .I1(n3750), .I2(n3744), .I3(n2967), 
            .O(n3751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5354.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5355 (.I0(\XI[15][25] ), .I1(\XI[14][25] ), .I2(n2954), 
            .I3(n2953), .O(n3752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5355.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5356 (.I0(\XI[13][25] ), .I1(\XI[12][25] ), .I2(n2953), 
            .I3(n2954), .O(n3753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5356.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5357 (.I0(n3752), .I1(n3753), .I2(n2959), .O(n3754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5357.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5358 (.I0(\XI[9][25] ), .I1(\XI[8][25] ), .I2(n2954), 
            .O(n3755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5358.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5359 (.I0(\XI[11][25] ), .I1(\XI[10][25] ), .I2(n2954), 
            .O(n3756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5359.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5360 (.I0(n3756), .I1(n3755), .I2(n2959), .I3(n2953), 
            .O(n3757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5360.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5361 (.I0(\XI[5][25] ), .I1(\XI[4][25] ), .I2(n2953), 
            .I3(n2954), .O(n3758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5361.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5362 (.I0(\XI[7][25] ), .I1(\XI[6][25] ), .I2(n2954), 
            .I3(n2953), .O(n3759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5362.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5366 (.I0(n3759), .I1(n3758), .I2(n3762), .I3(n2959), 
            .O(n3763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5366.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5367 (.I0(n3757), .I1(n3754), .I2(n3763), .I3(n2967), 
            .O(n3764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5367.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5368 (.I0(n3764), .I1(n3751), .I2(n3029), .I3(n2966), 
            .O(n3765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5368.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5369 (.I0(\PC[25] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5369.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5370 (.I0(n3764), .I1(n3751), .I2(n2991), .I3(n2966), 
            .O(n3767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5370.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5371 (.I0(n2983), .I1(\PC[25] ), .I2(n3383), .O(n3768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5371.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5372 (.I0(n3767), .I1(n3768), .I2(n3765), .I3(n3766), 
            .O(n501_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5372.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5373 (.I0(\XI[18][24] ), .I1(\XI[19][24] ), .I2(n51770), 
            .O(n3769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5373.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5374 (.I0(\XI[16][24] ), .I1(\XI[17][24] ), .I2(n51770), 
            .O(n3770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5374.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5375 (.I0(n3769), .I1(n3770), .I2(n2959), .I3(n2953), 
            .O(n3771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5375.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5376 (.I0(\XI[21][24] ), .I1(\XI[20][24] ), .I2(n2953), 
            .I3(n2954), .O(n3772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5376.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5377 (.I0(\XI[23][24] ), .I1(\XI[22][24] ), .I2(n51770), 
            .O(n3773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5377.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5378 (.I0(n3773), .I1(n3771), .I2(n3772), .I3(n2959), 
            .O(n3774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5378.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5379 (.I0(\XI[25][24] ), .I1(\XI[24][24] ), .I2(n2954), 
            .O(n3775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5379.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5380 (.I0(\XI[27][24] ), .I1(\XI[26][24] ), .I2(n2954), 
            .O(n3776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5380.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5381 (.I0(n3776), .I1(n3775), .I2(n2959), .I3(n2953), 
            .O(n3777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5381.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5382 (.I0(\XI[31][24] ), .I1(\XI[30][24] ), .I2(n2954), 
            .O(n3778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5382.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5383 (.I0(\XI[29][24] ), .I1(\XI[28][24] ), .I2(n2954), 
            .O(n3779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5383.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5384 (.I0(n3779), .I1(n3778), .I2(n2953), .I3(n2959), 
            .O(n3780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5384.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5385 (.I0(n3777), .I1(n3780), .I2(n3774), .I3(n2967), 
            .O(n3781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5385.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5386 (.I0(\XI[15][24] ), .I1(\XI[14][24] ), .I2(n2954), 
            .I3(n2953), .O(n3782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5386.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5387 (.I0(\XI[13][24] ), .I1(\XI[12][24] ), .I2(n2953), 
            .I3(n2954), .O(n3783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5387.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5388 (.I0(n3782), .I1(n3783), .I2(n2959), .O(n3784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5388.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5389 (.I0(\XI[9][24] ), .I1(\XI[8][24] ), .I2(n2954), 
            .O(n3785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5389.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5390 (.I0(\XI[11][24] ), .I1(\XI[10][24] ), .I2(n2954), 
            .O(n3786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5390.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5391 (.I0(n3786), .I1(n3785), .I2(n2959), .I3(n2953), 
            .O(n3787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5391.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5392 (.I0(\XI[5][24] ), .I1(\XI[4][24] ), .I2(n2953), 
            .I3(n2954), .O(n3788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5392.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5393 (.I0(\XI[7][24] ), .I1(\XI[6][24] ), .I2(n2954), 
            .I3(n2953), .O(n3789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5393.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5397 (.I0(n3789), .I1(n3788), .I2(n3792), .I3(n2959), 
            .O(n3793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5397.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5398 (.I0(n3787), .I1(n3784), .I2(n3793), .I3(n2967), 
            .O(n3794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5398.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5399 (.I0(n3794), .I1(n3781), .I2(n3029), .I3(n2966), 
            .O(n3795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5399.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5400 (.I0(\PC[24] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5400.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5401 (.I0(n3794), .I1(n3781), .I2(n2991), .I3(n2966), 
            .O(n3797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5401.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5402 (.I0(n2983), .I1(\PC[24] ), .I2(n3383), .O(n3798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5402.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5403 (.I0(n3797), .I1(n3798), .I2(n3795), .I3(n3796), 
            .O(n502_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5403.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5404 (.I0(\XI[18][31] ), .I1(\XI[19][31] ), .I2(n51770), 
            .O(n3799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5404.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5405 (.I0(\XI[16][31] ), .I1(\XI[17][31] ), .I2(n51770), 
            .O(n3800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5405.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5406 (.I0(n3799), .I1(n3800), .I2(n2959), .I3(n2953), 
            .O(n3801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5406.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5407 (.I0(\XI[21][31] ), .I1(\XI[20][31] ), .I2(n2953), 
            .I3(n2954), .O(n3802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5407.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5408 (.I0(\XI[23][31] ), .I1(\XI[22][31] ), .I2(n51770), 
            .O(n3803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5408.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5409 (.I0(n3803), .I1(n3801), .I2(n3802), .I3(n2959), 
            .O(n3804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5409.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5410 (.I0(\XI[25][31] ), .I1(\XI[24][31] ), .I2(n2954), 
            .O(n3805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5410.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5411 (.I0(\XI[27][31] ), .I1(\XI[26][31] ), .I2(n2954), 
            .O(n3806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5411.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5412 (.I0(n3806), .I1(n3805), .I2(n2959), .I3(n2953), 
            .O(n3807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5412.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5413 (.I0(\XI[31][31] ), .I1(\XI[30][31] ), .I2(n2954), 
            .O(n3808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5413.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5414 (.I0(\XI[29][31] ), .I1(\XI[28][31] ), .I2(n2954), 
            .O(n3809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5414.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5415 (.I0(n3809), .I1(n3808), .I2(n2953), .I3(n2959), 
            .O(n3810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5415.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5416 (.I0(n3807), .I1(n3810), .I2(n3804), .I3(n2967), 
            .O(n3811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5416.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5417 (.I0(\XI[15][31] ), .I1(\XI[14][31] ), .I2(n2954), 
            .I3(n2953), .O(n3812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5417.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5418 (.I0(\XI[13][31] ), .I1(\XI[12][31] ), .I2(n2953), 
            .I3(n2954), .O(n3813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5418.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5419 (.I0(n3812), .I1(n3813), .I2(n2959), .O(n3814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5419.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5420 (.I0(\XI[9][31] ), .I1(\XI[8][31] ), .I2(n2954), 
            .O(n3815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5420.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5421 (.I0(\XI[11][31] ), .I1(\XI[10][31] ), .I2(n2954), 
            .O(n3816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5421.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5422 (.I0(n3816), .I1(n3815), .I2(n2959), .I3(n2953), 
            .O(n3817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5422.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5423 (.I0(\XI[5][31] ), .I1(\XI[4][31] ), .I2(n2953), 
            .I3(n2954), .O(n3818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5423.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5424 (.I0(\XI[7][31] ), .I1(\XI[6][31] ), .I2(n2954), 
            .I3(n2953), .O(n3819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5424.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5428 (.I0(n3819), .I1(n3818), .I2(n3822), .I3(n2959), 
            .O(n3823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5428.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5429 (.I0(n3817), .I1(n3814), .I2(n3823), .I3(n2967), 
            .O(n3824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5429.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5430 (.I0(n3824), .I1(n3811), .I2(n3029), .I3(n2966), 
            .O(n3825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5430.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5431 (.I0(\PC[31] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5431.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5432 (.I0(n3824), .I1(n3811), .I2(n2991), .I3(n2966), 
            .O(n3827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5432.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5433 (.I0(n2983), .I1(\PC[31] ), .I2(n3383), .O(n3828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5433.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5434 (.I0(n3827), .I1(n3828), .I2(n3825), .I3(n3826), 
            .O(n495_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5434.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5435 (.I0(\XI[18][23] ), .I1(\XI[19][23] ), .I2(n51770), 
            .O(n3829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5435.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5436 (.I0(\XI[16][23] ), .I1(\XI[17][23] ), .I2(n51770), 
            .O(n3830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5436.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5437 (.I0(n3829), .I1(n3830), .I2(n2959), .I3(n2953), 
            .O(n3831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5437.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5438 (.I0(\XI[21][23] ), .I1(\XI[20][23] ), .I2(n2953), 
            .I3(n2954), .O(n3832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5438.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5439 (.I0(\XI[23][23] ), .I1(\XI[22][23] ), .I2(n51770), 
            .O(n3833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5439.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5440 (.I0(n3833), .I1(n3831), .I2(n3832), .I3(n2959), 
            .O(n3834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5440.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5441 (.I0(\XI[25][23] ), .I1(\XI[24][23] ), .I2(n2954), 
            .O(n3835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5441.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5442 (.I0(\XI[27][23] ), .I1(\XI[26][23] ), .I2(n2954), 
            .O(n3836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5442.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5443 (.I0(n3836), .I1(n3835), .I2(n2959), .I3(n2953), 
            .O(n3837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5443.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5444 (.I0(\XI[31][23] ), .I1(\XI[30][23] ), .I2(n2954), 
            .O(n3838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5444.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5445 (.I0(\XI[29][23] ), .I1(\XI[28][23] ), .I2(n2954), 
            .O(n3839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5445.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5446 (.I0(n3839), .I1(n3838), .I2(n2953), .I3(n2959), 
            .O(n3840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5446.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5447 (.I0(n3837), .I1(n3840), .I2(n3834), .I3(n2967), 
            .O(n3841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5447.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5448 (.I0(\XI[15][23] ), .I1(\XI[14][23] ), .I2(n2954), 
            .I3(n2953), .O(n3842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5448.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5449 (.I0(\XI[13][23] ), .I1(\XI[12][23] ), .I2(n2953), 
            .I3(n2954), .O(n3843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5449.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5450 (.I0(n3842), .I1(n3843), .I2(n2959), .O(n3844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5450.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5451 (.I0(\XI[9][23] ), .I1(\XI[8][23] ), .I2(n2954), 
            .O(n3845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5451.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5452 (.I0(\XI[11][23] ), .I1(\XI[10][23] ), .I2(n2954), 
            .O(n3846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5452.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5453 (.I0(n3846), .I1(n3845), .I2(n2959), .I3(n2953), 
            .O(n3847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5453.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5454 (.I0(\XI[5][23] ), .I1(\XI[4][23] ), .I2(n2953), 
            .I3(n2954), .O(n3848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5454.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5455 (.I0(\XI[7][23] ), .I1(\XI[6][23] ), .I2(n2954), 
            .I3(n2953), .O(n3849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5455.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5459 (.I0(n3849), .I1(n3848), .I2(n3852), .I3(n2959), 
            .O(n3853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5459.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5460 (.I0(n3847), .I1(n3844), .I2(n3853), .I3(n2967), 
            .O(n3854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5460.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5461 (.I0(n3854), .I1(n3841), .I2(n3029), .I3(n2966), 
            .O(n3855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5461.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5462 (.I0(\PC[23] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5462.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5463 (.I0(n3854), .I1(n3841), .I2(n2991), .I3(n2966), 
            .O(n3857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5463.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5464 (.I0(n2983), .I1(\PC[23] ), .I2(n3383), .O(n3858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5464.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5465 (.I0(n3857), .I1(n3858), .I2(n3855), .I3(n3856), 
            .O(n503_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5465.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5466 (.I0(\XI[18][30] ), .I1(\XI[19][30] ), .I2(n51770), 
            .O(n3859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5466.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5467 (.I0(\XI[16][30] ), .I1(\XI[17][30] ), .I2(n51770), 
            .O(n3860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5467.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5468 (.I0(n3859), .I1(n3860), .I2(n2959), .I3(n2953), 
            .O(n3861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5468.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5469 (.I0(\XI[21][30] ), .I1(\XI[20][30] ), .I2(n2953), 
            .I3(n2954), .O(n3862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5469.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5470 (.I0(\XI[23][30] ), .I1(\XI[22][30] ), .I2(n51770), 
            .O(n3863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5470.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5471 (.I0(n3863), .I1(n3861), .I2(n3862), .I3(n2959), 
            .O(n3864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5471.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5472 (.I0(\XI[25][30] ), .I1(\XI[24][30] ), .I2(n2954), 
            .O(n3865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5472.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5473 (.I0(\XI[27][30] ), .I1(\XI[26][30] ), .I2(n2954), 
            .O(n3866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5473.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5474 (.I0(n3866), .I1(n3865), .I2(n2959), .I3(n2953), 
            .O(n3867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5474.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5475 (.I0(\XI[31][30] ), .I1(\XI[30][30] ), .I2(n2954), 
            .O(n3868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5475.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5476 (.I0(\XI[29][30] ), .I1(\XI[28][30] ), .I2(n2954), 
            .O(n3869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5476.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5477 (.I0(n3869), .I1(n3868), .I2(n2953), .I3(n2959), 
            .O(n3870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5477.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5478 (.I0(n3867), .I1(n3870), .I2(n3864), .I3(n2967), 
            .O(n3871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5478.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5479 (.I0(\XI[15][30] ), .I1(\XI[14][30] ), .I2(n2954), 
            .I3(n2953), .O(n3872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5479.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5480 (.I0(\XI[13][30] ), .I1(\XI[12][30] ), .I2(n2953), 
            .I3(n2954), .O(n3873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5480.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5481 (.I0(n3872), .I1(n3873), .I2(n2959), .O(n3874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5481.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5482 (.I0(\XI[9][30] ), .I1(\XI[8][30] ), .I2(n2954), 
            .O(n3875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5482.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5483 (.I0(\XI[11][30] ), .I1(\XI[10][30] ), .I2(n2954), 
            .O(n3876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5483.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5484 (.I0(n3876), .I1(n3875), .I2(n2959), .I3(n2953), 
            .O(n3877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5484.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5485 (.I0(\XI[5][30] ), .I1(\XI[4][30] ), .I2(n2953), 
            .I3(n2954), .O(n3878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5485.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5486 (.I0(\XI[7][30] ), .I1(\XI[6][30] ), .I2(n2954), 
            .I3(n2953), .O(n3879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5486.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5490 (.I0(n3879), .I1(n3878), .I2(n3882), .I3(n2959), 
            .O(n3883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5490.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5491 (.I0(n3877), .I1(n3874), .I2(n3883), .I3(n2967), 
            .O(n3884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5491.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5492 (.I0(n3884), .I1(n3871), .I2(n3029), .I3(n2966), 
            .O(n3885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5492.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5493 (.I0(\PC[30] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5493.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5494 (.I0(n3884), .I1(n3871), .I2(n2991), .I3(n2966), 
            .O(n3887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5494.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5495 (.I0(n2983), .I1(\PC[30] ), .I2(n3383), .O(n3888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5495.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5496 (.I0(n3887), .I1(n3888), .I2(n3885), .I3(n3886), 
            .O(n496_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5496.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5497 (.I0(\XI[7][31] ), .I1(\XI[3][31] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n3889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5497.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5498 (.I0(\XI[5][31] ), .I1(\XI[1][31] ), .I2(n51786), 
            .I3(n3889), .O(n3890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5498.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5499 (.I0(\XI[6][31] ), .I1(\XI[2][31] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n3891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5499.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5500 (.I0(\XI[4][31] ), .I1(\XI[0][31] ), .I2(\INSTRUCTION[16] ), 
            .I3(n3891), .O(n3892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5500.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5501 (.I0(n3892), .I1(n3890), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n3893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5501.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5502 (.I0(\XI[11][31] ), .I1(\XI[9][31] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5502.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5503 (.I0(\XI[10][31] ), .I1(\XI[8][31] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5503.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5504 (.I0(\XI[15][31] ), .I1(\XI[13][31] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5504.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5505 (.I0(\XI[14][31] ), .I1(\XI[12][31] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5505.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5506 (.I0(n3897), .I1(n3896), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n3898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5506.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5507 (.I0(n3895), .I1(\INSTRUCTION[17] ), .I2(n3894), 
            .I3(n3898), .O(n3899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5507.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5508 (.I0(n3893), .I1(n3899), .I2(\INSTRUCTION[19] ), 
            .O(n3900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__5508.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__5509 (.I0(\XI[22][31] ), .I1(\XI[20][31] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n3901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5509.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5510 (.I0(\XI[18][31] ), .I1(\XI[16][31] ), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[16] ), .O(n3902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5510.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5511 (.I0(\XI[23][31] ), .I1(\XI[19][31] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n3903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5511.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5512 (.I0(\XI[21][31] ), .I1(\XI[17][31] ), .I2(n51786), 
            .I3(n3903), .O(n3904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5512.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5513 (.I0(n3902), .I1(n3901), .I2(n3904), .I3(\INSTRUCTION[15] ), 
            .O(n3905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__5513.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__5514 (.I0(\XI[27][31] ), .I1(\XI[25][31] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5514.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5515 (.I0(\XI[26][31] ), .I1(\XI[24][31] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5515.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5516 (.I0(\XI[31][31] ), .I1(\XI[29][31] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5516.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5517 (.I0(\XI[30][31] ), .I1(\XI[28][31] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5517.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5518 (.I0(n3909), .I1(n3908), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n3910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5518.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5519 (.I0(n3907), .I1(\INSTRUCTION[17] ), .I2(n3906), 
            .I3(n3910), .O(n3911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5519.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5520 (.I0(n3905), .I1(\INSTRUCTION[18] ), .I2(n3911), 
            .I3(\INSTRUCTION[19] ), .O(n3912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__5520.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__5521 (.I0(n2983), .I1(n51826), .I2(n3155), .O(n3913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__5521.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__5522 (.I0(n3912), .I1(n3900), .I2(n51726), .I3(n3913), 
            .O(n543_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5522.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5523 (.I0(\XI[18][22] ), .I1(\XI[19][22] ), .I2(n51770), 
            .O(n3914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5523.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5524 (.I0(\XI[16][22] ), .I1(\XI[17][22] ), .I2(n51770), 
            .O(n3915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__5524.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__5525 (.I0(n3914), .I1(n3915), .I2(n2959), .I3(n2953), 
            .O(n3916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5525.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5526 (.I0(\XI[21][22] ), .I1(\XI[20][22] ), .I2(n2953), 
            .I3(n2954), .O(n3917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5526.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5527 (.I0(\XI[23][22] ), .I1(\XI[22][22] ), .I2(n51770), 
            .O(n3918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5527.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5528 (.I0(n3918), .I1(n3916), .I2(n3917), .I3(n2959), 
            .O(n3919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e33 */ ;
    defparam LUT__5528.LUTMASK = 16'h0e33;
    EFX_LUT4 LUT__5529 (.I0(\XI[25][22] ), .I1(\XI[24][22] ), .I2(n2954), 
            .O(n3920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5529.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5530 (.I0(\XI[27][22] ), .I1(\XI[26][22] ), .I2(n2954), 
            .O(n3921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5530.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5531 (.I0(n3921), .I1(n3920), .I2(n2959), .I3(n2953), 
            .O(n3922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5531.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5532 (.I0(\XI[31][22] ), .I1(\XI[30][22] ), .I2(n2954), 
            .O(n3923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5532.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5533 (.I0(\XI[29][22] ), .I1(\XI[28][22] ), .I2(n2954), 
            .O(n3924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5533.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5534 (.I0(n3924), .I1(n3923), .I2(n2953), .I3(n2959), 
            .O(n3925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5534.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5535 (.I0(n3922), .I1(n3925), .I2(n3919), .I3(n2967), 
            .O(n3926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5535.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5536 (.I0(\XI[15][22] ), .I1(\XI[14][22] ), .I2(n2954), 
            .I3(n2953), .O(n3927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5536.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5537 (.I0(\XI[13][22] ), .I1(\XI[12][22] ), .I2(n2953), 
            .I3(n2954), .O(n3928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5537.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5538 (.I0(n3927), .I1(n3928), .I2(n2959), .O(n3929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5538.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5539 (.I0(\XI[9][22] ), .I1(\XI[8][22] ), .I2(n2954), 
            .O(n3930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5539.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5540 (.I0(\XI[11][22] ), .I1(\XI[10][22] ), .I2(n2954), 
            .O(n3931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5540.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5541 (.I0(n3931), .I1(n3930), .I2(n2959), .I3(n2953), 
            .O(n3932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5541.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5542 (.I0(\XI[5][22] ), .I1(\XI[4][22] ), .I2(n2953), 
            .I3(n2954), .O(n3933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5542.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5543 (.I0(\XI[7][22] ), .I1(\XI[6][22] ), .I2(n2954), 
            .I3(n2953), .O(n3934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5543.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5547 (.I0(n3934), .I1(n3933), .I2(n3937), .I3(n2959), 
            .O(n3938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5547.LUTMASK = 16'heef0;
    EFX_LUT4 \CutToMuxOpt_11/Lut_1  (.I0(\XI[0][13] ), .I1(\XI[1][13] ), 
            .I2(n2953), .I3(\CutToMuxOpt_11/n7 ), .O(n3438)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_11/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5548 (.I0(n3932), .I1(n3929), .I2(n3938), .I3(n2967), 
            .O(n3939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5548.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5549 (.I0(n3939), .I1(n3926), .I2(n3029), .I3(n2966), 
            .O(n3940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5549.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5550 (.I0(\PC[22] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5550.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5551 (.I0(n3939), .I1(n3926), .I2(n2991), .I3(n2966), 
            .O(n3942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__5551.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__5552 (.I0(n2983), .I1(\PC[22] ), .I2(n3383), .O(n3943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5552.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5553 (.I0(n3942), .I1(n3943), .I2(n3940), .I3(n3941), 
            .O(n504_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__5553.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__5554 (.I0(\XI[15][30] ), .I1(\XI[13][30] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5554.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5555 (.I0(\XI[14][30] ), .I1(\XI[12][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5555.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5556 (.I0(\XI[11][30] ), .I1(\XI[9][30] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5556.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5557 (.I0(\XI[10][30] ), .I1(\XI[8][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5557.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5558 (.I0(\XI[3][30] ), .I1(\XI[1][30] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5558.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5559 (.I0(n3946), .I1(n3947), .I2(n3948), .I3(\INSTRUCTION[18] ), 
            .O(n3949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5559.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5560 (.I0(n3944), .I1(n3945), .I2(n3949), .I3(\INSTRUCTION[17] ), 
            .O(n3950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5560.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5561 (.I0(\XI[6][30] ), .I1(\XI[4][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5561.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5562 (.I0(\XI[7][30] ), .I1(\XI[5][30] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5562.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5563 (.I0(\XI[2][30] ), .I1(\XI[0][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5563.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5564 (.I0(n3951), .I1(n3952), .I2(n3953), .I3(\INSTRUCTION[17] ), 
            .O(n3954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5564.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5565 (.I0(\INSTRUCTION[17] ), .I1(\INSTRUCTION[18] ), 
            .I2(n3954), .I3(n3950), .O(n3955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h03ce */ ;
    defparam LUT__5565.LUTMASK = 16'h03ce;
    EFX_LUT4 LUT__5566 (.I0(n2986), .I1(n51726), .I2(n3913), .O(n3956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__5566.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__5567 (.I0(n51730), .I1(n51826), .I2(n3956), .O(n3957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5567.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5568 (.I0(\XI[19][30] ), .I1(\XI[17][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5568.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5569 (.I0(\XI[16][30] ), .I1(\XI[18][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(n3958), .O(n3959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__5569.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__5570 (.I0(\XI[23][30] ), .I1(\XI[21][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5570.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5571 (.I0(\XI[22][30] ), .I1(\XI[20][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(n3960), .O(n3961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5571.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5572 (.I0(n3961), .I1(n3959), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n3962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5572.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5573 (.I0(\XI[31][30] ), .I1(\XI[29][30] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5573.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5574 (.I0(\XI[30][30] ), .I1(\XI[28][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5574.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5575 (.I0(\XI[27][30] ), .I1(\XI[25][30] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5575.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5576 (.I0(\XI[26][30] ), .I1(\XI[24][30] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5576.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5577 (.I0(\INSTRUCTION[17] ), .I1(n3966), .I2(n3965), 
            .I3(\INSTRUCTION[18] ), .O(n3967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5577.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5578 (.I0(n3964), .I1(n3963), .I2(\INSTRUCTION[17] ), 
            .I3(n3967), .O(n3968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5578.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5579 (.I0(n3962), .I1(n3968), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n3969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5579.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5580 (.I0(\INSTRUCTION[19] ), .I1(n3955), .I2(n3969), 
            .I3(n3957), .O(n544_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5580.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5581 (.I0(\XI[7][21] ), .I1(\XI[6][21] ), .I2(n2954), 
            .I3(n2953), .O(n3970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5581.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5582 (.I0(\XI[5][21] ), .I1(\XI[4][21] ), .I2(n2953), 
            .I3(n2954), .O(n3971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5582.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5583 (.I0(\XI[3][21] ), .I1(\XI[1][21] ), .I2(n2954), 
            .I3(n2953), .O(n3972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5583.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5584 (.I0(\XI[2][21] ), .I1(\XI[0][21] ), .I2(n2954), 
            .I3(n3972), .O(n3973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5584.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5585 (.I0(n3971), .I1(n3970), .I2(n3973), .I3(n2959), 
            .O(n3974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5585.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5586 (.I0(\XI[15][21] ), .I1(\XI[14][21] ), .I2(n2954), 
            .I3(n2953), .O(n3975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5586.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5587 (.I0(\XI[13][21] ), .I1(\XI[12][21] ), .I2(n2953), 
            .I3(n2954), .O(n3976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5587.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5588 (.I0(\XI[11][21] ), .I1(\XI[9][21] ), .I2(n2954), 
            .I3(n2953), .O(n3977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5588.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5589 (.I0(\XI[10][21] ), .I1(\XI[8][21] ), .I2(n2954), 
            .I3(n3977), .O(n3978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5589.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5590 (.I0(n3976), .I1(n3975), .I2(n3978), .I3(n2959), 
            .O(n3979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5590.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5591 (.I0(n3979), .I1(n3974), .I2(n2966), .I3(n2967), 
            .O(n3980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5591.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5592 (.I0(\XI[19][21] ), .I1(\XI[17][21] ), .I2(n2954), 
            .I3(n2953), .O(n3981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5592.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5593 (.I0(\XI[18][21] ), .I1(\XI[16][21] ), .I2(n2954), 
            .I3(n3981), .O(n3982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5593.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5594 (.I0(\XI[23][21] ), .I1(\XI[21][21] ), .I2(n2954), 
            .I3(n2953), .O(n3983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5594.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5595 (.I0(\XI[22][21] ), .I1(\XI[20][21] ), .I2(n2954), 
            .I3(n3983), .O(n3984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5595.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5596 (.I0(n3984), .I1(n3982), .I2(n2967), .I3(n2959), 
            .O(n3985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5596.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5597 (.I0(\XI[27][21] ), .I1(\XI[26][21] ), .I2(n2954), 
            .I3(n2953), .O(n3986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5597.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5598 (.I0(\XI[25][21] ), .I1(\XI[24][21] ), .I2(n2953), 
            .I3(n2954), .O(n3987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5598.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5599 (.I0(\XI[31][21] ), .I1(\XI[30][21] ), .I2(n2954), 
            .I3(n2953), .O(n3988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5599.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5600 (.I0(\XI[29][21] ), .I1(\XI[28][21] ), .I2(n2953), 
            .I3(n2954), .O(n3989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5600.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5601 (.I0(n3989), .I1(n3988), .I2(n2959), .I3(n2967), 
            .O(n3990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5601.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5602 (.I0(n3987), .I1(n2959), .I2(n3986), .I3(n3990), 
            .O(n3991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5602.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5603 (.I0(n3985), .I1(n3991), .I2(n2966), .O(n3992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5603.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5604 (.I0(n2983), .I1(\PC[21] ), .I2(n2986), .O(n3993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__5604.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__5605 (.I0(\PC[21] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n3994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__5605.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__5606 (.I0(n3994), .I1(n3029), .I2(n3993), .I3(n2991), 
            .O(n3995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__5606.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__5607 (.I0(n3992), .I1(n3980), .I2(n2987), .I3(n3995), 
            .O(n505_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__5607.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__5608 (.I0(\XI[3][29] ), .I1(\XI[1][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5608.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5609 (.I0(\XI[2][29] ), .I1(\XI[0][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(n3996), .O(n3997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5609.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5610 (.I0(\XI[6][29] ), .I1(\XI[4][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n3998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5610.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5611 (.I0(\XI[7][29] ), .I1(\XI[5][29] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n3999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5611.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5612 (.I0(n3999), .I1(n3998), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5612.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5613 (.I0(\INSTRUCTION[17] ), .I1(n3997), .I2(n4000), 
            .I3(\INSTRUCTION[19] ), .O(n4001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5613.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5614 (.I0(\INSTRUCTION[29] ), .I1(n51826), .I2(n3956), 
            .O(n4002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5614.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5615 (.I0(\XI[11][29] ), .I1(\XI[9][29] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5615.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5616 (.I0(\XI[10][29] ), .I1(\XI[8][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5616.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5617 (.I0(\XI[15][29] ), .I1(\XI[13][29] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5617.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5618 (.I0(\XI[14][29] ), .I1(\XI[12][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5618.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5619 (.I0(n4006), .I1(n4005), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5619.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5620 (.I0(n4004), .I1(\INSTRUCTION[17] ), .I2(n4003), 
            .I3(n4007), .O(n4008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5620.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5621 (.I0(\XI[19][29] ), .I1(\XI[17][29] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5621.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5622 (.I0(\XI[18][29] ), .I1(\XI[16][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5622.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5623 (.I0(\XI[23][29] ), .I1(\XI[21][29] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5623.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5624 (.I0(\XI[22][29] ), .I1(\XI[20][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5624.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5625 (.I0(n4012), .I1(n4011), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5625.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5626 (.I0(n4010), .I1(\INSTRUCTION[17] ), .I2(n4009), 
            .I3(n4013), .O(n4014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5626.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5627 (.I0(\XI[26][29] ), .I1(\XI[24][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5627.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5628 (.I0(\XI[27][29] ), .I1(\XI[25][29] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5628.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5629 (.I0(\XI[30][29] ), .I1(\XI[28][29] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5629.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5630 (.I0(\XI[31][29] ), .I1(\XI[29][29] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5630.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5631 (.I0(n4018), .I1(n4017), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5631.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5632 (.I0(n4016), .I1(\INSTRUCTION[17] ), .I2(n4015), 
            .I3(n4019), .O(n4020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5632.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5633 (.I0(n4020), .I1(n4014), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5633.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5634 (.I0(n4008), .I1(n4001), .I2(n4021), .I3(n4002), 
            .O(n545_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5634.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5635 (.I0(\XI[3][28] ), .I1(\XI[1][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5635.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5636 (.I0(\XI[2][28] ), .I1(\XI[0][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4022), .O(n4023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5636.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5637 (.I0(\XI[6][28] ), .I1(\XI[4][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5637.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5638 (.I0(\XI[7][28] ), .I1(\XI[5][28] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5638.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5639 (.I0(n4025), .I1(n4024), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5639.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5640 (.I0(\INSTRUCTION[17] ), .I1(n4023), .I2(n4026), 
            .I3(\INSTRUCTION[19] ), .O(n4027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5640.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5641 (.I0(\INSTRUCTION[28] ), .I1(n51826), .I2(n3956), 
            .O(n4028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5641.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5642 (.I0(\XI[11][28] ), .I1(\XI[9][28] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5642.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5643 (.I0(\XI[10][28] ), .I1(\XI[8][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5643.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5644 (.I0(\XI[15][28] ), .I1(\XI[13][28] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5644.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5645 (.I0(\XI[14][28] ), .I1(\XI[12][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5645.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5646 (.I0(n4032), .I1(n4031), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5646.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5647 (.I0(n4030), .I1(\INSTRUCTION[17] ), .I2(n4029), 
            .I3(n4033), .O(n4034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5647.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5648 (.I0(\XI[19][28] ), .I1(\XI[17][28] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5648.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5649 (.I0(\XI[18][28] ), .I1(\XI[16][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5649.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5650 (.I0(\XI[23][28] ), .I1(\XI[21][28] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5650.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5651 (.I0(\XI[22][28] ), .I1(\XI[20][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5651.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5652 (.I0(n4038), .I1(n4037), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5652.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5653 (.I0(n4036), .I1(\INSTRUCTION[17] ), .I2(n4035), 
            .I3(n4039), .O(n4040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5653.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5654 (.I0(\XI[26][28] ), .I1(\XI[24][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5654.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5655 (.I0(\XI[27][28] ), .I1(\XI[25][28] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5655.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5656 (.I0(\XI[30][28] ), .I1(\XI[28][28] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5656.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5657 (.I0(\XI[31][28] ), .I1(\XI[29][28] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5657.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5658 (.I0(n4044), .I1(n4043), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5658.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5659 (.I0(n4042), .I1(\INSTRUCTION[17] ), .I2(n4041), 
            .I3(n4045), .O(n4046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5659.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5660 (.I0(n4046), .I1(n4040), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5660.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5661 (.I0(n4034), .I1(n4027), .I2(n4047), .I3(n4028), 
            .O(n546_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5661.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5662 (.I0(\XI[3][27] ), .I1(\XI[1][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5662.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5663 (.I0(\XI[2][27] ), .I1(\XI[0][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4048), .O(n4049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5663.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5664 (.I0(\XI[6][27] ), .I1(\XI[4][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5664.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5665 (.I0(\XI[7][27] ), .I1(\XI[5][27] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5665.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5666 (.I0(n4051), .I1(n4050), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5666.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5667 (.I0(\INSTRUCTION[17] ), .I1(n4049), .I2(n4052), 
            .I3(\INSTRUCTION[19] ), .O(n4053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5667.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5668 (.I0(\INSTRUCTION[27] ), .I1(n51826), .I2(n3956), 
            .O(n4054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5668.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5669 (.I0(\XI[11][27] ), .I1(\XI[9][27] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5669.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5670 (.I0(\XI[10][27] ), .I1(\XI[8][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5670.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5671 (.I0(\XI[15][27] ), .I1(\XI[13][27] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5671.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5672 (.I0(\XI[14][27] ), .I1(\XI[12][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5672.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5673 (.I0(n4058), .I1(n4057), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5673.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5674 (.I0(n4056), .I1(\INSTRUCTION[17] ), .I2(n4055), 
            .I3(n4059), .O(n4060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5674.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5675 (.I0(\XI[19][27] ), .I1(\XI[17][27] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5675.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5676 (.I0(\XI[18][27] ), .I1(\XI[16][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5676.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5677 (.I0(\XI[23][27] ), .I1(\XI[21][27] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5677.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5678 (.I0(\XI[22][27] ), .I1(\XI[20][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5678.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5679 (.I0(n4064), .I1(n4063), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5679.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5680 (.I0(n4062), .I1(\INSTRUCTION[17] ), .I2(n4061), 
            .I3(n4065), .O(n4066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5680.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5681 (.I0(\XI[26][27] ), .I1(\XI[24][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5681.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5682 (.I0(\XI[27][27] ), .I1(\XI[25][27] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5682.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5683 (.I0(\XI[30][27] ), .I1(\XI[28][27] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5683.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5684 (.I0(\XI[31][27] ), .I1(\XI[29][27] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5684.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5685 (.I0(n4070), .I1(n4069), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5685.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5686 (.I0(n4068), .I1(\INSTRUCTION[17] ), .I2(n4067), 
            .I3(n4071), .O(n4072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5686.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5687 (.I0(n4072), .I1(n4066), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5687.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5688 (.I0(n4060), .I1(n4053), .I2(n4073), .I3(n4054), 
            .O(n547_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5688.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5689 (.I0(\XI[3][26] ), .I1(\XI[1][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5689.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5690 (.I0(\XI[2][26] ), .I1(\XI[0][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4074), .O(n4075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5690.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5691 (.I0(\XI[6][26] ), .I1(\XI[4][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5691.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5692 (.I0(\XI[7][26] ), .I1(\XI[5][26] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5692.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5693 (.I0(n4077), .I1(n4076), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5693.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5694 (.I0(\INSTRUCTION[17] ), .I1(n4075), .I2(n4078), 
            .I3(\INSTRUCTION[19] ), .O(n4079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5694.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5695 (.I0(\INSTRUCTION[26] ), .I1(n51826), .I2(n3956), 
            .O(n4080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5695.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5696 (.I0(\XI[11][26] ), .I1(\XI[9][26] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5696.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5697 (.I0(\XI[10][26] ), .I1(\XI[8][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5697.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5698 (.I0(\XI[15][26] ), .I1(\XI[13][26] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5698.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5699 (.I0(\XI[14][26] ), .I1(\XI[12][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5699.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5700 (.I0(n4084), .I1(n4083), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5700.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5701 (.I0(n4082), .I1(\INSTRUCTION[17] ), .I2(n4081), 
            .I3(n4085), .O(n4086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5701.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5702 (.I0(\XI[19][26] ), .I1(\XI[17][26] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5702.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5703 (.I0(\XI[18][26] ), .I1(\XI[16][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5703.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5704 (.I0(\XI[23][26] ), .I1(\XI[21][26] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5704.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5705 (.I0(\XI[22][26] ), .I1(\XI[20][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5705.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5706 (.I0(n4090), .I1(n4089), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5706.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5707 (.I0(n4088), .I1(\INSTRUCTION[17] ), .I2(n4087), 
            .I3(n4091), .O(n4092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5707.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5708 (.I0(\XI[26][26] ), .I1(\XI[24][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5708.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5709 (.I0(\XI[27][26] ), .I1(\XI[25][26] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5709.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5710 (.I0(\XI[30][26] ), .I1(\XI[28][26] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5710.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5711 (.I0(\XI[31][26] ), .I1(\XI[29][26] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5711.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5712 (.I0(n4096), .I1(n4095), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5712.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5713 (.I0(n4094), .I1(\INSTRUCTION[17] ), .I2(n4093), 
            .I3(n4097), .O(n4098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5713.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5714 (.I0(n4098), .I1(n4092), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5714.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5715 (.I0(n4086), .I1(n4079), .I2(n4099), .I3(n4080), 
            .O(n548_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5715.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5716 (.I0(\XI[3][25] ), .I1(\XI[1][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5716.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5717 (.I0(\XI[2][25] ), .I1(\XI[0][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4100), .O(n4101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5717.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5718 (.I0(\XI[6][25] ), .I1(\XI[4][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5718.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5719 (.I0(\XI[7][25] ), .I1(\XI[5][25] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5719.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5720 (.I0(n4103), .I1(n4102), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5720.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5721 (.I0(\INSTRUCTION[17] ), .I1(n4101), .I2(n4104), 
            .I3(\INSTRUCTION[19] ), .O(n4105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5721.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5722 (.I0(\INSTRUCTION[25] ), .I1(n51826), .I2(n3956), 
            .O(n4106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5722.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5723 (.I0(\XI[11][25] ), .I1(\XI[9][25] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5723.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5724 (.I0(\XI[10][25] ), .I1(\XI[8][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5724.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5725 (.I0(\XI[15][25] ), .I1(\XI[13][25] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5725.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5726 (.I0(\XI[14][25] ), .I1(\XI[12][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5726.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5727 (.I0(n4110), .I1(n4109), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5727.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5728 (.I0(n4108), .I1(\INSTRUCTION[17] ), .I2(n4107), 
            .I3(n4111), .O(n4112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5728.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5729 (.I0(\XI[19][25] ), .I1(\XI[17][25] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5729.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5730 (.I0(\XI[18][25] ), .I1(\XI[16][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5730.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5731 (.I0(\XI[23][25] ), .I1(\XI[21][25] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5731.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5732 (.I0(\XI[22][25] ), .I1(\XI[20][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5732.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5733 (.I0(n4116), .I1(n4115), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5733.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5734 (.I0(n4114), .I1(\INSTRUCTION[17] ), .I2(n4113), 
            .I3(n4117), .O(n4118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5734.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5735 (.I0(\XI[26][25] ), .I1(\XI[24][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5735.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5736 (.I0(\XI[27][25] ), .I1(\XI[25][25] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5736.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5737 (.I0(\XI[30][25] ), .I1(\XI[28][25] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5737.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5738 (.I0(\XI[31][25] ), .I1(\XI[29][25] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5738.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5739 (.I0(n4122), .I1(n4121), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5739.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5740 (.I0(n4120), .I1(\INSTRUCTION[17] ), .I2(n4119), 
            .I3(n4123), .O(n4124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5740.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5741 (.I0(n4124), .I1(n4118), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5741.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5742 (.I0(n4112), .I1(n4105), .I2(n4125), .I3(n4106), 
            .O(n549_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5742.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5743 (.I0(\XI[3][24] ), .I1(\XI[1][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5743.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5744 (.I0(\XI[2][24] ), .I1(\XI[0][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4126), .O(n4127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5744.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5745 (.I0(\XI[6][24] ), .I1(\XI[4][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5745.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5746 (.I0(\XI[7][24] ), .I1(\XI[5][24] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5746.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5747 (.I0(n4129), .I1(n4128), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5747.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5748 (.I0(\INSTRUCTION[17] ), .I1(n4127), .I2(n4130), 
            .I3(\INSTRUCTION[19] ), .O(n4131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5748.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5749 (.I0(n2966), .I1(n51826), .I2(n3956), .O(n4132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5749.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5750 (.I0(\XI[11][24] ), .I1(\XI[9][24] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5750.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5751 (.I0(\XI[10][24] ), .I1(\XI[8][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5751.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5752 (.I0(\XI[15][24] ), .I1(\XI[13][24] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5752.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5753 (.I0(\XI[14][24] ), .I1(\XI[12][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5753.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5754 (.I0(n4136), .I1(n4135), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5754.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5755 (.I0(n4134), .I1(\INSTRUCTION[17] ), .I2(n4133), 
            .I3(n4137), .O(n4138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5755.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5756 (.I0(\XI[19][24] ), .I1(\XI[17][24] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5756.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5757 (.I0(\XI[18][24] ), .I1(\XI[16][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5757.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5758 (.I0(\XI[23][24] ), .I1(\XI[21][24] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5758.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5759 (.I0(\XI[22][24] ), .I1(\XI[20][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5759.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5760 (.I0(n4142), .I1(n4141), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5760.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5761 (.I0(n4140), .I1(\INSTRUCTION[17] ), .I2(n4139), 
            .I3(n4143), .O(n4144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5761.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5762 (.I0(\XI[26][24] ), .I1(\XI[24][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5762.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5763 (.I0(\XI[27][24] ), .I1(\XI[25][24] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5763.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5764 (.I0(\XI[30][24] ), .I1(\XI[28][24] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5764.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5765 (.I0(\XI[31][24] ), .I1(\XI[29][24] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5765.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5766 (.I0(n4148), .I1(n4147), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5766.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5767 (.I0(n4146), .I1(\INSTRUCTION[17] ), .I2(n4145), 
            .I3(n4149), .O(n4150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5767.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5768 (.I0(n4150), .I1(n4144), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5768.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5769 (.I0(n4138), .I1(n4131), .I2(n4151), .I3(n4132), 
            .O(n550_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5769.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5770 (.I0(\XI[3][23] ), .I1(\XI[1][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5770.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5771 (.I0(\XI[2][23] ), .I1(\XI[0][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4152), .O(n4153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5771.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5772 (.I0(\XI[6][23] ), .I1(\XI[4][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5772.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5773 (.I0(\XI[7][23] ), .I1(\XI[5][23] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5773.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5774 (.I0(n4155), .I1(n4154), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5774.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5775 (.I0(\INSTRUCTION[17] ), .I1(n4153), .I2(n4156), 
            .I3(\INSTRUCTION[19] ), .O(n4157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5775.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5776 (.I0(n2967), .I1(n51826), .I2(n3956), .O(n4158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5776.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5777 (.I0(\XI[11][23] ), .I1(\XI[9][23] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5777.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5778 (.I0(\XI[10][23] ), .I1(\XI[8][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5778.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5779 (.I0(\XI[15][23] ), .I1(\XI[13][23] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5779.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5780 (.I0(\XI[14][23] ), .I1(\XI[12][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5780.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5781 (.I0(n4162), .I1(n4161), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5781.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5782 (.I0(n4160), .I1(\INSTRUCTION[17] ), .I2(n4159), 
            .I3(n4163), .O(n4164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5782.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5783 (.I0(\XI[19][23] ), .I1(\XI[17][23] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5783.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5784 (.I0(\XI[18][23] ), .I1(\XI[16][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5784.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5785 (.I0(\XI[23][23] ), .I1(\XI[21][23] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5785.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5786 (.I0(\XI[22][23] ), .I1(\XI[20][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5786.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5787 (.I0(n4168), .I1(n4167), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5787.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5788 (.I0(n4166), .I1(\INSTRUCTION[17] ), .I2(n4165), 
            .I3(n4169), .O(n4170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5788.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5789 (.I0(\XI[26][23] ), .I1(\XI[24][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5789.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5790 (.I0(\XI[27][23] ), .I1(\XI[25][23] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5790.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5791 (.I0(\XI[30][23] ), .I1(\XI[28][23] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5791.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5792 (.I0(\XI[31][23] ), .I1(\XI[29][23] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5792.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5793 (.I0(n4174), .I1(n4173), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5793.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5794 (.I0(n4172), .I1(\INSTRUCTION[17] ), .I2(n4171), 
            .I3(n4175), .O(n4176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5794.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5795 (.I0(n4176), .I1(n4170), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5795.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5796 (.I0(n4164), .I1(n4157), .I2(n4177), .I3(n4158), 
            .O(n551_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5796.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5797 (.I0(\XI[3][22] ), .I1(\XI[1][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5797.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5798 (.I0(\XI[2][22] ), .I1(\XI[0][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4178), .O(n4179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5798.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5799 (.I0(\XI[6][22] ), .I1(\XI[4][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5799.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5800 (.I0(\XI[7][22] ), .I1(\XI[5][22] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5800.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5801 (.I0(n4181), .I1(n4180), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5801.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5802 (.I0(\INSTRUCTION[17] ), .I1(n4179), .I2(n4182), 
            .I3(\INSTRUCTION[19] ), .O(n4183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5802.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5803 (.I0(n2959), .I1(n51826), .I2(n3956), .O(n4184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5803.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5804 (.I0(\XI[11][22] ), .I1(\XI[9][22] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5804.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5805 (.I0(\XI[10][22] ), .I1(\XI[8][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5805.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5806 (.I0(\XI[15][22] ), .I1(\XI[13][22] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5806.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5807 (.I0(\XI[14][22] ), .I1(\XI[12][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5807.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5808 (.I0(n4188), .I1(n4187), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5808.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5809 (.I0(n4186), .I1(\INSTRUCTION[17] ), .I2(n4185), 
            .I3(n4189), .O(n4190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5809.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5810 (.I0(\XI[19][22] ), .I1(\XI[17][22] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5810.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5811 (.I0(\XI[18][22] ), .I1(\XI[16][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5811.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5812 (.I0(\XI[23][22] ), .I1(\XI[21][22] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5812.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5813 (.I0(\XI[22][22] ), .I1(\XI[20][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5813.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5814 (.I0(n4194), .I1(n4193), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5814.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5815 (.I0(n4192), .I1(\INSTRUCTION[17] ), .I2(n4191), 
            .I3(n4195), .O(n4196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5815.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5816 (.I0(\XI[26][22] ), .I1(\XI[24][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5816.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5817 (.I0(\XI[27][22] ), .I1(\XI[25][22] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5817.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5818 (.I0(\XI[30][22] ), .I1(\XI[28][22] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5818.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5819 (.I0(\XI[31][22] ), .I1(\XI[29][22] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5819.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5820 (.I0(n4200), .I1(n4199), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5820.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5821 (.I0(n4198), .I1(\INSTRUCTION[17] ), .I2(n4197), 
            .I3(n4201), .O(n4202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5821.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5822 (.I0(n4202), .I1(n4196), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5822.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5823 (.I0(n4190), .I1(n4183), .I2(n4203), .I3(n4184), 
            .O(n552_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5823.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5824 (.I0(\XI[3][21] ), .I1(\XI[1][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5824.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5825 (.I0(\XI[2][21] ), .I1(\XI[0][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4204), .O(n4205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5825.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5826 (.I0(\XI[6][21] ), .I1(\XI[4][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5826.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5827 (.I0(\XI[7][21] ), .I1(\XI[5][21] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5827.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5828 (.I0(n4207), .I1(n4206), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5828.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5829 (.I0(\INSTRUCTION[17] ), .I1(n4205), .I2(n4208), 
            .I3(\INSTRUCTION[19] ), .O(n4209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5829.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5830 (.I0(n2953), .I1(n51826), .I2(n3956), .O(n4210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5830.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5831 (.I0(\XI[11][21] ), .I1(\XI[9][21] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5831.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5832 (.I0(\XI[10][21] ), .I1(\XI[8][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5832.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5833 (.I0(\XI[15][21] ), .I1(\XI[13][21] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5833.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5834 (.I0(\XI[14][21] ), .I1(\XI[12][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5834.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5835 (.I0(n4214), .I1(n4213), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5835.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5836 (.I0(n4212), .I1(\INSTRUCTION[17] ), .I2(n4211), 
            .I3(n4215), .O(n4216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5836.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5837 (.I0(\XI[19][21] ), .I1(\XI[17][21] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5837.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5838 (.I0(\XI[18][21] ), .I1(\XI[16][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5838.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5839 (.I0(\XI[23][21] ), .I1(\XI[21][21] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5839.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5840 (.I0(\XI[22][21] ), .I1(\XI[20][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5840.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5841 (.I0(n4220), .I1(n4219), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5841.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5842 (.I0(n4218), .I1(\INSTRUCTION[17] ), .I2(n4217), 
            .I3(n4221), .O(n4222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5842.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5843 (.I0(\XI[26][21] ), .I1(\XI[24][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5843.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5844 (.I0(\XI[27][21] ), .I1(\XI[25][21] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5844.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5845 (.I0(\XI[30][21] ), .I1(\XI[28][21] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5845.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5846 (.I0(\XI[31][21] ), .I1(\XI[29][21] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5846.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5847 (.I0(n4226), .I1(n4225), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5847.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5848 (.I0(n4224), .I1(\INSTRUCTION[17] ), .I2(n4223), 
            .I3(n4227), .O(n4228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5848.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5849 (.I0(n4228), .I1(n4222), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5849.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5850 (.I0(n4216), .I1(n4209), .I2(n4229), .I3(n4210), 
            .O(n553_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5850.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5851 (.I0(\XI[26][20] ), .I1(\XI[24][20] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5851.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5852 (.I0(\XI[27][20] ), .I1(\XI[25][20] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5852.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5853 (.I0(\XI[30][20] ), .I1(\XI[28][20] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5853.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5854 (.I0(\XI[31][20] ), .I1(\XI[29][20] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5854.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5855 (.I0(n4233), .I1(n4232), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5855.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5856 (.I0(n4231), .I1(\INSTRUCTION[17] ), .I2(n4230), 
            .I3(n4234), .O(n4235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5856.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5857 (.I0(\XI[19][20] ), .I1(\XI[17][20] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5857.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5858 (.I0(\XI[18][20] ), .I1(\XI[16][20] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5858.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5859 (.I0(\XI[23][20] ), .I1(\XI[21][20] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5859.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5860 (.I0(\XI[22][20] ), .I1(\XI[20][20] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5860.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5861 (.I0(n4239), .I1(n4238), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5861.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5862 (.I0(n4237), .I1(\INSTRUCTION[17] ), .I2(n4236), 
            .I3(n4240), .O(n4241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5862.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5863 (.I0(n4235), .I1(n4241), .I2(\INSTRUCTION[19] ), 
            .O(n4242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5863.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5864 (.I0(\XI[7][20] ), .I1(\XI[5][20] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5864.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5865 (.I0(\XI[6][20] ), .I1(\XI[4][20] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5865.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5866 (.I0(n4244), .I1(n4243), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5866.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5867 (.I0(\XI[2][20] ), .I1(\XI[0][20] ), .I2(\INSTRUCTION[16] ), 
            .O(n4246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5867.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5868 (.I0(\XI[3][20] ), .I1(\XI[1][20] ), .I2(\INSTRUCTION[16] ), 
            .O(n4247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5868.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5869 (.I0(n4247), .I1(n4246), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[15] ), .O(n4248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5869.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5870 (.I0(\XI[10][20] ), .I1(\XI[8][20] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5870.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5871 (.I0(\XI[11][20] ), .I1(\XI[9][20] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5871.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5872 (.I0(\XI[14][20] ), .I1(\XI[12][20] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5872.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5873 (.I0(\XI[15][20] ), .I1(\XI[13][20] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5873.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5874 (.I0(n4252), .I1(n4251), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5874.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5875 (.I0(n4250), .I1(\INSTRUCTION[17] ), .I2(n4249), 
            .I3(n4253), .O(n4254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5875.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5876 (.I0(n4248), .I1(n4245), .I2(n4254), .I3(\INSTRUCTION[19] ), 
            .O(n4255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__5876.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__5877 (.I0(n2954), .I1(n51826), .I2(n3956), .O(n4256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5877.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5878 (.I0(n4255), .I1(n4242), .I2(n3913), .I3(n4256), 
            .O(n554_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5878.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5879 (.I0(\XI[3][19] ), .I1(\XI[1][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5879.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5880 (.I0(\XI[2][19] ), .I1(\XI[0][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4257), .O(n4258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5880.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5881 (.I0(\XI[10][19] ), .I1(\XI[8][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5881.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5882 (.I0(\XI[11][19] ), .I1(\XI[9][19] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5882.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5883 (.I0(n4260), .I1(n4259), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5883.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5884 (.I0(\INSTRUCTION[18] ), .I1(n4258), .I2(n4261), 
            .I3(\INSTRUCTION[19] ), .O(n4262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__5884.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__5885 (.I0(\INSTRUCTION[19] ), .I1(n51826), .I2(n3956), 
            .O(n4263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__5885.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__5886 (.I0(\XI[7][19] ), .I1(\XI[5][19] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5886.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5887 (.I0(\XI[6][19] ), .I1(\XI[4][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5887.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5888 (.I0(\XI[15][19] ), .I1(\XI[13][19] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5888.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5889 (.I0(\XI[14][19] ), .I1(\XI[12][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5889.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5890 (.I0(n4267), .I1(n4266), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5890.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5891 (.I0(n4265), .I1(\INSTRUCTION[18] ), .I2(n4264), 
            .I3(n4268), .O(n4269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5891.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5892 (.I0(\XI[19][19] ), .I1(\XI[17][19] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5892.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5893 (.I0(\XI[18][19] ), .I1(\XI[16][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5893.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5894 (.I0(\XI[27][19] ), .I1(\XI[25][19] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5894.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5895 (.I0(\XI[26][19] ), .I1(\XI[24][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5895.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5896 (.I0(n4273), .I1(n4272), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5896.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5897 (.I0(n4271), .I1(\INSTRUCTION[18] ), .I2(n4270), 
            .I3(n4274), .O(n4275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5897.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5898 (.I0(\XI[22][19] ), .I1(\XI[20][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5898.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5899 (.I0(\XI[23][19] ), .I1(\XI[21][19] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5899.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5900 (.I0(\XI[30][19] ), .I1(\XI[28][19] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5900.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5901 (.I0(\XI[31][19] ), .I1(\XI[29][19] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5901.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5902 (.I0(n4279), .I1(n4278), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5902.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5903 (.I0(n4277), .I1(\INSTRUCTION[18] ), .I2(n4276), 
            .I3(n4280), .O(n4281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5903.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5904 (.I0(n4281), .I1(n4275), .I2(\INSTRUCTION[19] ), 
            .I3(n3913), .O(n4282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5904.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5905 (.I0(n4269), .I1(n4262), .I2(n4282), .I3(n4263), 
            .O(n555_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__5905.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__5906 (.I0(\INSTRUCTION[19] ), .I1(\INSTRUCTION[18] ), 
            .I2(n3174), .O(n4283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__5906.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__5907 (.I0(\XI[7][18] ), .I1(\XI[5][18] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5907.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5908 (.I0(\XI[6][18] ), .I1(\XI[4][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5908.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5909 (.I0(\XI[15][18] ), .I1(\XI[13][18] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5909.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5910 (.I0(\XI[14][18] ), .I1(\XI[12][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5910.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5911 (.I0(n4287), .I1(n4286), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5911.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5912 (.I0(n4285), .I1(\INSTRUCTION[18] ), .I2(n4284), 
            .I3(n4288), .O(n4289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5912.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5913 (.I0(\XI[3][18] ), .I1(\XI[1][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5913.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5914 (.I0(\XI[0][18] ), .I1(\XI[2][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4290), .O(n4291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__5914.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__5915 (.I0(\XI[11][18] ), .I1(\XI[9][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5915.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5916 (.I0(\XI[10][18] ), .I1(\XI[8][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4292), .O(n4293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5916.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5917 (.I0(n4293), .I1(n4291), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__5917.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__5918 (.I0(n3155), .I1(n4289), .I2(n4294), .O(n4295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__5918.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__5919 (.I0(\XI[30][18] ), .I1(\XI[28][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5919.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5920 (.I0(\XI[31][18] ), .I1(\XI[29][18] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5920.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5921 (.I0(\XI[23][18] ), .I1(\XI[21][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5921.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5922 (.I0(\XI[22][18] ), .I1(\XI[20][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4298), .O(n4299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5922.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5923 (.I0(n4296), .I1(n4297), .I2(n4299), .I3(\INSTRUCTION[18] ), 
            .O(n4300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__5923.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__5924 (.I0(\XI[19][18] ), .I1(\XI[17][18] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5924.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5925 (.I0(\XI[18][18] ), .I1(\XI[16][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5925.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5926 (.I0(\XI[27][18] ), .I1(\XI[25][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5926.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5927 (.I0(\XI[26][18] ), .I1(\XI[24][18] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4303), .O(n4304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5927.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5928 (.I0(n4302), .I1(n4301), .I2(n4304), .I3(\INSTRUCTION[18] ), 
            .O(n4305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__5928.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__5929 (.I0(n4305), .I1(n4300), .I2(n3155), .I3(\INSTRUCTION[17] ), 
            .O(n4306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5929.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5930 (.I0(n4295), .I1(n4306), .I2(n3174), .I3(n4283), 
            .O(n556_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0af3 */ ;
    defparam LUT__5930.LUTMASK = 16'h0af3;
    EFX_LUT4 LUT__5931 (.I0(\INSTRUCTION[17] ), .I1(\INSTRUCTION[18] ), 
            .I2(n51826), .I3(n3913), .O(n4307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__5931.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__5932 (.I0(\XI[22][17] ), .I1(\XI[18][17] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5932.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5933 (.I0(\XI[20][17] ), .I1(\XI[16][17] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4308), .O(n4309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5933.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5934 (.I0(\XI[23][17] ), .I1(\XI[19][17] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5934.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5935 (.I0(\XI[21][17] ), .I1(\XI[17][17] ), .I2(n51786), 
            .I3(n4310), .O(n4311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5935.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5936 (.I0(n4311), .I1(n4309), .I2(\INSTRUCTION[19] ), 
            .I3(\INSTRUCTION[15] ), .O(n4312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__5936.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__5937 (.I0(\XI[6][17] ), .I1(\XI[2][17] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5937.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5938 (.I0(\XI[4][17] ), .I1(\XI[0][17] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4313), .O(n4314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5938.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5939 (.I0(\XI[7][17] ), .I1(\XI[3][17] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5939.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5940 (.I0(\XI[5][17] ), .I1(\XI[1][17] ), .I2(n51786), 
            .I3(n4315), .O(n4316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5940.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5941 (.I0(n4316), .I1(n4314), .I2(\INSTRUCTION[19] ), 
            .I3(n4312), .O(n4317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__5941.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__5942 (.I0(\XI[27][17] ), .I1(\XI[25][17] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5942.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5943 (.I0(\XI[26][17] ), .I1(\XI[24][17] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5943.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5944 (.I0(\XI[31][17] ), .I1(\XI[29][17] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5944.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5945 (.I0(\XI[30][17] ), .I1(\XI[28][17] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5945.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5946 (.I0(n4321), .I1(n4320), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5946.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5947 (.I0(n4319), .I1(\INSTRUCTION[17] ), .I2(n4318), 
            .I3(n4322), .O(n4323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5947.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5948 (.I0(\XI[11][17] ), .I1(\XI[9][17] ), .I2(\INSTRUCTION[16] ), 
            .O(n4324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5948.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5949 (.I0(\XI[10][17] ), .I1(\XI[8][17] ), .I2(\INSTRUCTION[16] ), 
            .O(n4325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5949.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5950 (.I0(n4325), .I1(n4324), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[15] ), .O(n4326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__5950.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__5951 (.I0(\XI[15][17] ), .I1(\XI[13][17] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5951.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5952 (.I0(\XI[14][17] ), .I1(\XI[12][17] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5952.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5953 (.I0(n4328), .I1(n4327), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5953.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5954 (.I0(n4326), .I1(n4329), .I2(n4323), .I3(\INSTRUCTION[19] ), 
            .O(n4330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__5954.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__5955 (.I0(n4317), .I1(n4307), .I2(n4330), .I3(n3913), 
            .O(n557_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7033 */ ;
    defparam LUT__5955.LUTMASK = 16'h7033;
    EFX_LUT4 LUT__5956 (.I0(\XI[15][16] ), .I1(\XI[13][16] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5956.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5957 (.I0(\XI[14][16] ), .I1(\XI[12][16] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5957.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5958 (.I0(n4332), .I1(n4331), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5958.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5959 (.I0(\XI[11][16] ), .I1(\XI[9][16] ), .I2(\INSTRUCTION[16] ), 
            .O(n4334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5959.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5960 (.I0(\XI[10][16] ), .I1(\XI[8][16] ), .I2(\INSTRUCTION[16] ), 
            .O(n4335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5960.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5961 (.I0(n4335), .I1(n4334), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[15] ), .O(n4336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__5961.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__5962 (.I0(\XI[7][16] ), .I1(\XI[3][16] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5962.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5963 (.I0(\XI[5][16] ), .I1(\XI[1][16] ), .I2(n51786), 
            .I3(n4337), .O(n4338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5963.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5964 (.I0(\XI[6][16] ), .I1(\XI[2][16] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5964.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5965 (.I0(\XI[4][16] ), .I1(\XI[0][16] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4339), .O(n4340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5965.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5966 (.I0(n4340), .I1(n4338), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5966.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5967 (.I0(n4336), .I1(n4333), .I2(n4341), .I3(\INSTRUCTION[19] ), 
            .O(n4342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__5967.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__5968 (.I0(\XI[23][16] ), .I1(\XI[19][16] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5968.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5969 (.I0(\XI[21][16] ), .I1(\XI[17][16] ), .I2(n51786), 
            .I3(n4343), .O(n4344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5969.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5970 (.I0(\XI[22][16] ), .I1(\XI[18][16] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5970.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5971 (.I0(\XI[20][16] ), .I1(\XI[16][16] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4345), .O(n4346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5971.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5972 (.I0(n4346), .I1(n4344), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5972.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5973 (.I0(\XI[27][16] ), .I1(\XI[25][16] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5973.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5974 (.I0(\XI[26][16] ), .I1(\XI[24][16] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5974.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5975 (.I0(\XI[31][16] ), .I1(\XI[29][16] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5975.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5976 (.I0(\XI[30][16] ), .I1(\XI[28][16] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5976.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5977 (.I0(n4351), .I1(n4350), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__5977.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__5978 (.I0(n4349), .I1(\INSTRUCTION[17] ), .I2(n4348), 
            .I3(n4352), .O(n4353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__5978.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__5979 (.I0(n4347), .I1(n4353), .I2(\INSTRUCTION[19] ), 
            .O(n4354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5979.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5980 (.I0(\INSTRUCTION[17] ), .I1(\INSTRUCTION[16] ), 
            .I2(n51826), .O(n4355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5980.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5981 (.I0(n4354), .I1(n4342), .I2(n4355), .I3(n3913), 
            .O(n558_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__5981.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__5982 (.I0(\XI[2][15] ), .I1(\XI[0][15] ), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[16] ), .O(n4356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5982.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5983 (.I0(\XI[6][15] ), .I1(\XI[4][15] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5983.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5984 (.I0(\XI[7][15] ), .I1(\XI[3][15] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__5984.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__5985 (.I0(\XI[5][15] ), .I1(\XI[1][15] ), .I2(n51786), 
            .I3(n4358), .O(n4359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__5985.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__5986 (.I0(n4357), .I1(n4356), .I2(n4359), .I3(\INSTRUCTION[15] ), 
            .O(n4360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__5986.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__5987 (.I0(\XI[14][15] ), .I1(\XI[12][15] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5987.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5988 (.I0(\XI[15][15] ), .I1(\XI[13][15] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5988.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__5989 (.I0(\XI[10][15] ), .I1(\XI[8][15] ), .I2(\INSTRUCTION[16] ), 
            .O(n4363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5989.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5990 (.I0(\XI[11][15] ), .I1(\XI[9][15] ), .I2(\INSTRUCTION[16] ), 
            .O(n4364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5990.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5991 (.I0(n4364), .I1(n4363), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[15] ), .O(n4365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5991.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5992 (.I0(n4362), .I1(n4361), .I2(\INSTRUCTION[17] ), 
            .I3(n4365), .O(n4366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__5992.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__5993 (.I0(n4366), .I1(n4360), .I2(\INSTRUCTION[19] ), 
            .I3(\INSTRUCTION[18] ), .O(n4367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__5993.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__5994 (.I0(\XI[23][15] ), .I1(\XI[19][15] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5994.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5995 (.I0(\XI[21][15] ), .I1(\XI[17][15] ), .I2(n51786), 
            .I3(n4368), .O(n4369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5995.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5996 (.I0(\XI[22][15] ), .I1(\XI[18][15] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__5996.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__5997 (.I0(\XI[20][15] ), .I1(\XI[16][15] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4370), .O(n4371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__5997.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__5998 (.I0(n4371), .I1(n4369), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5998.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5999 (.I0(\XI[27][15] ), .I1(\XI[25][15] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__5999.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6000 (.I0(\XI[26][15] ), .I1(\XI[24][15] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6000.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6001 (.I0(\XI[31][15] ), .I1(\XI[29][15] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6001.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6002 (.I0(\XI[30][15] ), .I1(\XI[28][15] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6002.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6003 (.I0(n4376), .I1(n4375), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6003.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6004 (.I0(n4374), .I1(\INSTRUCTION[17] ), .I2(n4373), 
            .I3(n4377), .O(n4378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6004.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6005 (.I0(n4372), .I1(n4378), .I2(\INSTRUCTION[19] ), 
            .O(n4379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6005.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6006 (.I0(\INSTRUCTION[15] ), .I1(\INSTRUCTION[16] ), 
            .I2(n51826), .O(n4380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6006.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6007 (.I0(n4379), .I1(n4367), .I2(n4380), .I3(n3913), 
            .O(n559_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__6007.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__6008 (.I0(n51794), .I1(n51790), .I2(n51826), .O(n4381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6008.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6009 (.I0(\XI[7][14] ), .I1(\XI[3][14] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6009.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6010 (.I0(\XI[1][14] ), .I1(\XI[5][14] ), .I2(n51786), 
            .I3(n4382), .O(n4383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__6010.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__6011 (.I0(\XI[6][14] ), .I1(\XI[2][14] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6011.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6012 (.I0(\XI[4][14] ), .I1(\XI[0][14] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4384), .O(n4385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6012.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6013 (.I0(n4385), .I1(n4383), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__6013.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__6014 (.I0(\XI[27][14] ), .I1(\XI[25][14] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6014.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6015 (.I0(\XI[26][14] ), .I1(\XI[24][14] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6015.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6016 (.I0(\XI[31][14] ), .I1(\XI[29][14] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6016.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6017 (.I0(\XI[30][14] ), .I1(\XI[28][14] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6017.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6018 (.I0(n4390), .I1(n4389), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6018.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6019 (.I0(n4388), .I1(\INSTRUCTION[17] ), .I2(n4387), 
            .I3(n4391), .O(n4392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6019.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6020 (.I0(\XI[17][14] ), .I1(\XI[19][14] ), .I2(n51786), 
            .O(n4393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6020.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6021 (.I0(\XI[21][14] ), .I1(\XI[23][14] ), .I2(n51786), 
            .O(n4394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6021.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6022 (.I0(n4394), .I1(n4393), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[15] ), .O(n4395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6022.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6023 (.I0(\XI[22][14] ), .I1(\XI[20][14] ), .I2(\INSTRUCTION[16] ), 
            .O(n4396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6023.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6024 (.I0(\XI[18][14] ), .I1(\XI[16][14] ), .I2(\INSTRUCTION[16] ), 
            .O(n4397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6024.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6025 (.I0(n4397), .I1(n4396), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[17] ), .O(n4398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6025.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6026 (.I0(n4398), .I1(\INSTRUCTION[18] ), .I2(n4395), 
            .I3(\INSTRUCTION[19] ), .O(n4399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6026.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6027 (.I0(\XI[11][14] ), .I1(\XI[9][14] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6027.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6028 (.I0(\XI[10][14] ), .I1(\XI[8][14] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4400), .O(n4401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6028.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6029 (.I0(\XI[15][14] ), .I1(\XI[13][14] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6029.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6030 (.I0(\XI[14][14] ), .I1(\XI[12][14] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6030.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6031 (.I0(n4403), .I1(n4402), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6031.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6032 (.I0(\INSTRUCTION[17] ), .I1(n4401), .I2(n4404), 
            .I3(\INSTRUCTION[19] ), .O(n4405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6032.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6033 (.I0(n4392), .I1(n4399), .I2(n4386), .I3(n4405), 
            .O(n4406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6033.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6034 (.I0(n4406), .I1(n4381), .I2(n3913), .O(n560_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6034.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6035 (.I0(\XI[7][13] ), .I1(\XI[3][13] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6035.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6036 (.I0(\XI[5][13] ), .I1(\XI[1][13] ), .I2(n51786), 
            .I3(n4407), .O(n4408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6036.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6037 (.I0(\XI[6][13] ), .I1(\XI[2][13] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6037.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6038 (.I0(\XI[4][13] ), .I1(\XI[0][13] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4409), .O(n4410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6038.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6039 (.I0(n4410), .I1(n4408), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6039.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6040 (.I0(\XI[11][13] ), .I1(\XI[9][13] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6040.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6041 (.I0(\XI[10][13] ), .I1(\XI[8][13] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6041.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6042 (.I0(\XI[15][13] ), .I1(\XI[13][13] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6042.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6043 (.I0(\XI[14][13] ), .I1(\XI[12][13] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6043.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6044 (.I0(n4415), .I1(n4414), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6044.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6045 (.I0(n4413), .I1(\INSTRUCTION[17] ), .I2(n4412), 
            .I3(n4416), .O(n4417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6045.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6046 (.I0(n4411), .I1(n4417), .I2(\INSTRUCTION[19] ), 
            .O(n4418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6046.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6047 (.I0(\XI[22][13] ), .I1(\XI[20][13] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6047.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6048 (.I0(\XI[18][13] ), .I1(\XI[16][13] ), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[16] ), .O(n4420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6048.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6049 (.I0(\XI[23][13] ), .I1(\XI[19][13] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6049.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6050 (.I0(\XI[21][13] ), .I1(\XI[17][13] ), .I2(n51786), 
            .I3(n4421), .O(n4422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6050.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6051 (.I0(n4420), .I1(n4419), .I2(n4422), .I3(\INSTRUCTION[15] ), 
            .O(n4423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6051.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6052 (.I0(\XI[27][13] ), .I1(\XI[25][13] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6052.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6053 (.I0(\XI[26][13] ), .I1(\XI[24][13] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6053.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6054 (.I0(\XI[31][13] ), .I1(\XI[29][13] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6054.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6055 (.I0(\XI[30][13] ), .I1(\XI[28][13] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6055.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6056 (.I0(n4427), .I1(n4426), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6056.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6057 (.I0(n4425), .I1(\INSTRUCTION[17] ), .I2(n4424), 
            .I3(n4428), .O(n4429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6057.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6058 (.I0(n4423), .I1(\INSTRUCTION[18] ), .I2(n4429), 
            .I3(\INSTRUCTION[19] ), .O(n4430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6058.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6059 (.I0(n51794), .I1(n51798), .I2(n51826), .O(n4431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6059.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6060 (.I0(n4430), .I1(n4418), .I2(n4431), .I3(n3913), 
            .O(n561_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__6060.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__6061 (.I0(\XI[14][12] ), .I1(\XI[12][12] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6061.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6062 (.I0(\XI[15][12] ), .I1(\XI[13][12] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6062.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6063 (.I0(\XI[11][12] ), .I1(\XI[9][12] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6063.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6064 (.I0(\XI[10][12] ), .I1(\XI[8][12] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4434), .O(n4435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6064.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6065 (.I0(n4432), .I1(n4433), .I2(n4435), .I3(\INSTRUCTION[17] ), 
            .O(n4436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6065.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6066 (.I0(\XI[6][12] ), .I1(\XI[4][12] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6066.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6067 (.I0(\XI[2][12] ), .I1(\XI[0][12] ), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[16] ), .O(n4438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6067.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6068 (.I0(\XI[7][12] ), .I1(\XI[3][12] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6068.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6069 (.I0(\XI[5][12] ), .I1(\XI[1][12] ), .I2(n51786), 
            .I3(n4439), .O(n4440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6069.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6070 (.I0(n4438), .I1(n4437), .I2(n4440), .I3(\INSTRUCTION[15] ), 
            .O(n4441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6070.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6071 (.I0(n4441), .I1(n4436), .I2(\INSTRUCTION[19] ), 
            .I3(\INSTRUCTION[18] ), .O(n4442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6071.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6072 (.I0(\XI[23][12] ), .I1(\XI[19][12] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6072.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6073 (.I0(\XI[21][12] ), .I1(\XI[17][12] ), .I2(n51786), 
            .I3(n4443), .O(n4444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6073.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6074 (.I0(\XI[22][12] ), .I1(\XI[18][12] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6074.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6075 (.I0(\XI[20][12] ), .I1(\XI[16][12] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4445), .O(n4446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6075.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6076 (.I0(n4446), .I1(n4444), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6076.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6077 (.I0(\XI[27][12] ), .I1(\XI[25][12] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6077.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6078 (.I0(\XI[26][12] ), .I1(\XI[24][12] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6078.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6079 (.I0(\XI[31][12] ), .I1(\XI[29][12] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6079.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6080 (.I0(\XI[30][12] ), .I1(\XI[28][12] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6080.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6081 (.I0(n4451), .I1(n4450), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6081.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6082 (.I0(n4449), .I1(\INSTRUCTION[17] ), .I2(n4448), 
            .I3(n4452), .O(n4453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6082.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6083 (.I0(n4447), .I1(n4453), .I2(\INSTRUCTION[19] ), 
            .O(n4454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6083.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6084 (.I0(n51802), .I1(n51798), .I2(n51826), .O(n4455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6084.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6085 (.I0(n4454), .I1(n4442), .I2(n4455), .I3(n3913), 
            .O(n562_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__6085.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__6086 (.I0(\XI[3][11] ), .I1(\XI[1][11] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6086.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6087 (.I0(\XI[0][11] ), .I1(\XI[2][11] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4456), .O(n4457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__6087.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__6088 (.I0(\XI[7][11] ), .I1(\XI[5][11] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6088.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6089 (.I0(\XI[6][11] ), .I1(\XI[4][11] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4458), .O(n4459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6089.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6090 (.I0(n4459), .I1(n4457), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__6090.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__6091 (.I0(\XI[15][11] ), .I1(\XI[13][11] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6091.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6092 (.I0(\XI[14][11] ), .I1(\XI[12][11] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6092.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6093 (.I0(\XI[11][11] ), .I1(\XI[9][11] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6093.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6094 (.I0(\XI[10][11] ), .I1(\XI[8][11] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6094.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6095 (.I0(\INSTRUCTION[17] ), .I1(n4464), .I2(n4463), 
            .I3(\INSTRUCTION[18] ), .O(n4465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6095.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6096 (.I0(n4462), .I1(n4461), .I2(\INSTRUCTION[17] ), 
            .I3(n4465), .O(n4466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6096.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6097 (.I0(\INSTRUCTION[19] ), .I1(n4460), .I2(n4466), 
            .I3(n3155), .O(n4467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__6097.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__6098 (.I0(\XI[18][11] ), .I1(\XI[16][11] ), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[16] ), .O(n4468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6098.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6099 (.I0(\XI[26][11] ), .I1(\XI[24][11] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[18] ), .O(n4469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6099.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6100 (.I0(\XI[27][11] ), .I1(\XI[19][11] ), .I2(n51786), 
            .I3(\INSTRUCTION[18] ), .O(n4470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__6100.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__6101 (.I0(\XI[25][11] ), .I1(\XI[17][11] ), .I2(n51786), 
            .I3(n4470), .O(n4471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__6101.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__6102 (.I0(n4469), .I1(n4468), .I2(n4471), .I3(\INSTRUCTION[15] ), 
            .O(n4472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6102.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6103 (.I0(\XI[30][11] ), .I1(\XI[28][11] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6103.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6104 (.I0(\XI[31][11] ), .I1(\XI[29][11] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6104.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6105 (.I0(\XI[22][11] ), .I1(\XI[20][11] ), .I2(\INSTRUCTION[16] ), 
            .O(n4475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6105.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6106 (.I0(\XI[23][11] ), .I1(\XI[21][11] ), .I2(\INSTRUCTION[16] ), 
            .O(n4476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6106.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6107 (.I0(n4476), .I1(n4475), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6107.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6108 (.I0(n4474), .I1(n4473), .I2(\INSTRUCTION[18] ), 
            .I3(n4477), .O(n4478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6108.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6109 (.I0(n4478), .I1(n4472), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[19] ), .O(n4479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6109.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6110 (.I0(n3155), .I1(n51802), .I2(n3174), .O(n4480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6110.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6111 (.I0(n4479), .I1(n4467), .I2(n4480), .O(n563_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6111.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6112 (.I0(\XI[15][10] ), .I1(\XI[13][10] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6112.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6113 (.I0(\XI[14][10] ), .I1(\XI[12][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6113.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6114 (.I0(\XI[11][10] ), .I1(\XI[9][10] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6114.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6115 (.I0(\XI[10][10] ), .I1(\XI[8][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6115.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6116 (.I0(\INSTRUCTION[17] ), .I1(n4484), .I2(n4483), 
            .I3(\INSTRUCTION[18] ), .O(n4485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6116.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6117 (.I0(n4482), .I1(n4481), .I2(\INSTRUCTION[17] ), 
            .I3(n4485), .O(n4486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6117.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6118 (.I0(\INSTRUCTION[19] ), .I1(n4486), .I2(n51770), 
            .I3(n3155), .O(n4487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__6118.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__6119 (.I0(\XI[31][10] ), .I1(\XI[29][10] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6119.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6120 (.I0(\XI[30][10] ), .I1(\XI[28][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6120.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6121 (.I0(\XI[23][10] ), .I1(\XI[21][10] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6121.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6122 (.I0(\XI[22][10] ), .I1(\XI[20][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6122.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6123 (.I0(n4491), .I1(\INSTRUCTION[18] ), .I2(n4490), 
            .I3(\INSTRUCTION[17] ), .O(n4492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6123.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6124 (.I0(n4489), .I1(n4488), .I2(\INSTRUCTION[18] ), 
            .I3(n4492), .O(n4493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6124.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6125 (.I0(\XI[7][10] ), .I1(\XI[3][10] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6125.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6126 (.I0(\XI[5][10] ), .I1(\XI[1][10] ), .I2(n51786), 
            .I3(n4494), .O(n4495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6126.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6127 (.I0(\XI[6][10] ), .I1(\XI[2][10] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6127.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6128 (.I0(\XI[4][10] ), .I1(\XI[0][10] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4496), .O(n4497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6128.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6129 (.I0(n4497), .I1(n4495), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6129.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6130 (.I0(\XI[19][10] ), .I1(\XI[17][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6130.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6131 (.I0(\XI[18][10] ), .I1(\XI[16][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4499), .O(n4500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6131.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6132 (.I0(\XI[27][10] ), .I1(\XI[25][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6132.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6133 (.I0(\XI[26][10] ), .I1(\XI[24][10] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4501), .O(n4502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6133.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6134 (.I0(n4502), .I1(n4500), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6134.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6135 (.I0(n4493), .I1(n4503), .I2(n4498), .I3(\INSTRUCTION[19] ), 
            .O(n4504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6135.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6136 (.I0(n4504), .I1(n3155), .I2(n3174), .I3(n4487), 
            .O(n564_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6136.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6137 (.I0(\XI[15][9] ), .I1(\XI[13][9] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6137.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6138 (.I0(\XI[14][9] ), .I1(\XI[12][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6138.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6139 (.I0(\XI[11][9] ), .I1(\XI[9][9] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6139.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6140 (.I0(\XI[10][9] ), .I1(\XI[8][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6140.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6141 (.I0(\INSTRUCTION[17] ), .I1(n4508), .I2(n4507), 
            .I3(\INSTRUCTION[18] ), .O(n4509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6141.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6142 (.I0(n4506), .I1(n4505), .I2(\INSTRUCTION[17] ), 
            .I3(n4509), .O(n4510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6142.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6143 (.I0(\INSTRUCTION[19] ), .I1(n4510), .I2(n51730), 
            .I3(n3155), .O(n4511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__6143.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__6144 (.I0(\XI[31][9] ), .I1(\XI[29][9] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6144.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6145 (.I0(\XI[30][9] ), .I1(\XI[28][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6145.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6146 (.I0(\XI[23][9] ), .I1(\XI[21][9] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6146.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6147 (.I0(\XI[22][9] ), .I1(\XI[20][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6147.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6148 (.I0(n4515), .I1(\INSTRUCTION[18] ), .I2(n4514), 
            .I3(\INSTRUCTION[17] ), .O(n4516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6148.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6149 (.I0(n4513), .I1(n4512), .I2(\INSTRUCTION[18] ), 
            .I3(n4516), .O(n4517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6149.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6150 (.I0(\XI[7][9] ), .I1(\XI[3][9] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6150.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6151 (.I0(\XI[5][9] ), .I1(\XI[1][9] ), .I2(n51786), 
            .I3(n4518), .O(n4519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6151.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6152 (.I0(\XI[6][9] ), .I1(\XI[2][9] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6152.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6153 (.I0(\XI[4][9] ), .I1(\XI[0][9] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4520), .O(n4521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6153.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6154 (.I0(n4521), .I1(n4519), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6154.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6155 (.I0(\XI[19][9] ), .I1(\XI[17][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6155.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6156 (.I0(\XI[18][9] ), .I1(\XI[16][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4523), .O(n4524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6156.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6157 (.I0(\XI[27][9] ), .I1(\XI[25][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6157.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6158 (.I0(\XI[26][9] ), .I1(\XI[24][9] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4525), .O(n4526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6158.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6159 (.I0(n4526), .I1(n4524), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6159.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6160 (.I0(n4517), .I1(n4527), .I2(n4522), .I3(\INSTRUCTION[19] ), 
            .O(n4528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6160.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6161 (.I0(n4528), .I1(n3155), .I2(n3174), .I3(n4511), 
            .O(n565_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6161.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6162 (.I0(\XI[3][8] ), .I1(\XI[1][8] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6162.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6163 (.I0(\XI[0][8] ), .I1(\XI[2][8] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4529), .O(n4530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__6163.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__6164 (.I0(\XI[7][8] ), .I1(\XI[5][8] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6164.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6165 (.I0(\XI[6][8] ), .I1(\XI[4][8] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4531), .O(n4532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6165.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6166 (.I0(n4532), .I1(n4530), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__6166.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__6167 (.I0(\XI[15][8] ), .I1(\XI[13][8] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6167.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6168 (.I0(\XI[14][8] ), .I1(\XI[12][8] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6168.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6169 (.I0(\XI[11][8] ), .I1(\XI[9][8] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6169.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6170 (.I0(\XI[10][8] ), .I1(\XI[8][8] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6170.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6171 (.I0(\INSTRUCTION[17] ), .I1(n4537), .I2(n4536), 
            .I3(\INSTRUCTION[18] ), .O(n4538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6171.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6172 (.I0(n4535), .I1(n4534), .I2(\INSTRUCTION[17] ), 
            .I3(n4538), .O(n4539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6172.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6173 (.I0(\INSTRUCTION[19] ), .I1(n4533), .I2(n4539), 
            .I3(n3155), .O(n4540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__6173.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__6174 (.I0(\XI[18][8] ), .I1(\XI[16][8] ), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[16] ), .O(n4541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6174.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6175 (.I0(\XI[26][8] ), .I1(\XI[24][8] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[18] ), .O(n4542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6175.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6176 (.I0(\XI[27][8] ), .I1(\XI[19][8] ), .I2(n51786), 
            .I3(\INSTRUCTION[18] ), .O(n4543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6176.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6177 (.I0(\XI[25][8] ), .I1(\XI[17][8] ), .I2(n51786), 
            .I3(n4543), .O(n4544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6177.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6178 (.I0(n4542), .I1(n4541), .I2(n4544), .I3(\INSTRUCTION[15] ), 
            .O(n4545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6178.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6179 (.I0(\XI[30][8] ), .I1(\XI[28][8] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6179.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6180 (.I0(\XI[31][8] ), .I1(\XI[29][8] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6180.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6181 (.I0(\XI[22][8] ), .I1(\XI[20][8] ), .I2(\INSTRUCTION[16] ), 
            .O(n4548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6181.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6182 (.I0(\XI[23][8] ), .I1(\XI[21][8] ), .I2(\INSTRUCTION[16] ), 
            .O(n4549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6182.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6183 (.I0(n4549), .I1(n4548), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6183.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6184 (.I0(n4547), .I1(n4546), .I2(\INSTRUCTION[18] ), 
            .I3(n4550), .O(n4551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6184.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6185 (.I0(n4551), .I1(n4545), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[19] ), .O(n4552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6185.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6186 (.I0(n3155), .I1(n51734), .I2(n3174), .O(n4553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6186.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6187 (.I0(n4552), .I1(n4540), .I2(n4553), .O(n566_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6187.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6188 (.I0(\XII[15][7] ), .I1(\XII[13][7] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6188.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6189 (.I0(\XII[14][7] ), .I1(\XII[12][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6189.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6190 (.I0(\XII[11][7] ), .I1(\XII[9][7] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6190.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6191 (.I0(\XII[10][7] ), .I1(\XII[8][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6191.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6192 (.I0(\INSTRUCTION[17] ), .I1(n4557), .I2(n4556), 
            .I3(\INSTRUCTION[18] ), .O(n4558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6192.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6193 (.I0(n4555), .I1(n4554), .I2(\INSTRUCTION[17] ), 
            .I3(n4558), .O(n4559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6193.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6194 (.I0(\INSTRUCTION[19] ), .I1(n4559), .I2(n51738), 
            .I3(n3155), .O(n4560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__6194.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__6195 (.I0(\XII[31][7] ), .I1(\XII[29][7] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6195.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6196 (.I0(\XII[30][7] ), .I1(\XII[28][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6196.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6197 (.I0(\XII[23][7] ), .I1(\XII[21][7] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6197.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6198 (.I0(\XII[22][7] ), .I1(\XII[20][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6198.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6199 (.I0(n4564), .I1(\INSTRUCTION[18] ), .I2(n4563), 
            .I3(\INSTRUCTION[17] ), .O(n4565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6199.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6200 (.I0(n4562), .I1(n4561), .I2(\INSTRUCTION[18] ), 
            .I3(n4565), .O(n4566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6200.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6201 (.I0(\XII[7][7] ), .I1(\XII[3][7] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6201.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6202 (.I0(\XII[5][7] ), .I1(\XII[1][7] ), .I2(n51786), 
            .I3(n4567), .O(n4568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6202.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6203 (.I0(\XII[6][7] ), .I1(\XII[2][7] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6203.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6204 (.I0(\XII[4][7] ), .I1(\XII[0][7] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4569), .O(n4570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6204.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6205 (.I0(n4570), .I1(n4568), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6205.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6206 (.I0(\XII[19][7] ), .I1(\XII[17][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6206.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6207 (.I0(\XII[18][7] ), .I1(\XII[16][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4572), .O(n4573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6207.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6208 (.I0(\XII[27][7] ), .I1(\XII[25][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6208.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6209 (.I0(\XII[26][7] ), .I1(\XII[24][7] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4574), .O(n4575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6209.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6210 (.I0(n4575), .I1(n4573), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6210.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6211 (.I0(n4566), .I1(n4576), .I2(n4571), .I3(\INSTRUCTION[19] ), 
            .O(n4577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6211.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6212 (.I0(n4577), .I1(n3155), .I2(n3174), .I3(n4560), 
            .O(n567_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6212.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6213 (.I0(\XII[15][6] ), .I1(\XII[13][6] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6213.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6214 (.I0(\XII[14][6] ), .I1(\XII[12][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6214.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6215 (.I0(\XII[11][6] ), .I1(\XII[9][6] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6215.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6216 (.I0(\XII[10][6] ), .I1(\XII[8][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6216.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6217 (.I0(\INSTRUCTION[17] ), .I1(n4581), .I2(n4580), 
            .I3(\INSTRUCTION[18] ), .O(n4582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6217.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6218 (.I0(n4579), .I1(n4578), .I2(\INSTRUCTION[17] ), 
            .I3(n4582), .O(n4583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6218.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6219 (.I0(\INSTRUCTION[19] ), .I1(n4583), .I2(n51742), 
            .I3(n3155), .O(n4584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__6219.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__6220 (.I0(\XII[31][6] ), .I1(\XII[29][6] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6220.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6221 (.I0(\XII[30][6] ), .I1(\XII[28][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6221.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6222 (.I0(\XII[23][6] ), .I1(\XII[21][6] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6222.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6223 (.I0(\XII[22][6] ), .I1(\XII[20][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6223.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6224 (.I0(n4588), .I1(\INSTRUCTION[18] ), .I2(n4587), 
            .I3(\INSTRUCTION[17] ), .O(n4589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6224.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6225 (.I0(n4586), .I1(n4585), .I2(\INSTRUCTION[18] ), 
            .I3(n4589), .O(n4590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6225.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6226 (.I0(\XII[7][6] ), .I1(\XII[3][6] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6226.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6227 (.I0(\XII[5][6] ), .I1(\XII[1][6] ), .I2(n51786), 
            .I3(n4591), .O(n4592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6227.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6228 (.I0(\XII[6][6] ), .I1(\XII[2][6] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6228.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6229 (.I0(\XII[4][6] ), .I1(\XII[0][6] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4593), .O(n4594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6229.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6230 (.I0(n4594), .I1(n4592), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6230.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6231 (.I0(\XII[19][6] ), .I1(\XII[17][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6231.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6232 (.I0(\XII[18][6] ), .I1(\XII[16][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4596), .O(n4597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6232.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6233 (.I0(\XII[27][6] ), .I1(\XII[25][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6233.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6234 (.I0(\XII[26][6] ), .I1(\XII[24][6] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4598), .O(n4599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6234.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6235 (.I0(n4599), .I1(n4597), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6235.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6236 (.I0(n4590), .I1(n4600), .I2(n4595), .I3(\INSTRUCTION[19] ), 
            .O(n4601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6236.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6237 (.I0(n4601), .I1(n3155), .I2(n3174), .I3(n4584), 
            .O(n568_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6237.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6238 (.I0(\XII[15][5] ), .I1(\XII[13][5] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6238.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6239 (.I0(\XII[14][5] ), .I1(\XII[12][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6239.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6240 (.I0(\XII[11][5] ), .I1(\XII[9][5] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6240.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6241 (.I0(\XII[10][5] ), .I1(\XII[8][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6241.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6242 (.I0(\INSTRUCTION[17] ), .I1(n4605), .I2(n4604), 
            .I3(\INSTRUCTION[18] ), .O(n4606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6242.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6243 (.I0(n4603), .I1(n4602), .I2(\INSTRUCTION[17] ), 
            .I3(n4606), .O(n4607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6243.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6244 (.I0(\INSTRUCTION[19] ), .I1(n4607), .I2(n51746), 
            .I3(n3155), .O(n4608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__6244.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__6245 (.I0(\XII[31][5] ), .I1(\XII[29][5] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6245.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6246 (.I0(\XII[30][5] ), .I1(\XII[28][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6246.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6247 (.I0(\XII[23][5] ), .I1(\XII[21][5] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6247.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6248 (.I0(\XII[22][5] ), .I1(\XII[20][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6248.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6249 (.I0(n4612), .I1(\INSTRUCTION[18] ), .I2(n4611), 
            .I3(\INSTRUCTION[17] ), .O(n4613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6249.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6250 (.I0(n4610), .I1(n4609), .I2(\INSTRUCTION[18] ), 
            .I3(n4613), .O(n4614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6250.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6251 (.I0(\XII[7][5] ), .I1(\XII[3][5] ), .I2(n51786), 
            .I3(\INSTRUCTION[17] ), .O(n4615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6251.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6252 (.I0(\XII[5][5] ), .I1(\XII[1][5] ), .I2(n51786), 
            .I3(n4615), .O(n4616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6252.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6253 (.I0(\XII[6][5] ), .I1(\XII[2][5] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[17] ), .O(n4617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6253.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6254 (.I0(\XII[4][5] ), .I1(\XII[0][5] ), .I2(\INSTRUCTION[16] ), 
            .I3(n4617), .O(n4618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6254.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6255 (.I0(n4618), .I1(n4616), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6255.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6256 (.I0(\XII[19][5] ), .I1(\XII[17][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6256.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6257 (.I0(\XII[18][5] ), .I1(\XII[16][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4620), .O(n4621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6257.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6258 (.I0(\XII[27][5] ), .I1(\XII[25][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6258.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6259 (.I0(\XII[26][5] ), .I1(\XII[24][5] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4622), .O(n4623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6259.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6260 (.I0(n4623), .I1(n4621), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[18] ), .O(n4624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6260.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6261 (.I0(n4614), .I1(n4624), .I2(n4619), .I3(\INSTRUCTION[19] ), 
            .O(n4625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6261.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6262 (.I0(n4625), .I1(n3155), .I2(n3174), .I3(n4608), 
            .O(n569_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6262.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6263 (.I0(\XII[26][4] ), .I1(\XII[24][4] ), .I2(\INSTRUCTION[16] ), 
            .O(n4626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6263.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6264 (.I0(\XII[18][4] ), .I1(\XII[16][4] ), .I2(\INSTRUCTION[16] ), 
            .O(n4627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6264.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6265 (.I0(n4627), .I1(n4626), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[18] ), .O(n4628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6265.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6266 (.I0(\XII[17][4] ), .I1(\XII[19][4] ), .I2(n51786), 
            .O(n4629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6266.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6267 (.I0(\XII[25][4] ), .I1(\XII[27][4] ), .I2(n51786), 
            .O(n4630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6267.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6268 (.I0(n4630), .I1(n4629), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6268.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6269 (.I0(\XII[22][4] ), .I1(\XII[20][4] ), .I2(\INSTRUCTION[16] ), 
            .O(n4632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6269.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6270 (.I0(\XII[23][4] ), .I1(\XII[21][4] ), .I2(\INSTRUCTION[16] ), 
            .O(n4633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6270.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6271 (.I0(n4633), .I1(n4632), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6271.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6272 (.I0(\XII[30][4] ), .I1(\XII[28][4] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6272.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6273 (.I0(\XII[31][4] ), .I1(\XII[29][4] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6273.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6274 (.I0(n4635), .I1(n4636), .I2(\INSTRUCTION[18] ), 
            .O(n4637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6274.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6275 (.I0(n4637), .I1(n4634), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[19] ), .O(n4638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6275.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6276 (.I0(n4631), .I1(\INSTRUCTION[17] ), .I2(n4628), 
            .I3(n4638), .O(n4639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6276.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6277 (.I0(\XII[3][4] ), .I1(\XII[1][4] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6277.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6278 (.I0(\XII[2][4] ), .I1(\XII[0][4] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4640), .O(n4641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6278.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6279 (.I0(\XII[7][4] ), .I1(\XII[5][4] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6279.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6280 (.I0(\XII[6][4] ), .I1(\XII[4][4] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4642), .O(n4643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6280.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6281 (.I0(n4643), .I1(n4641), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6281.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6282 (.I0(\XII[15][4] ), .I1(\XII[13][4] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6282.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6283 (.I0(\XII[14][4] ), .I1(\XII[12][4] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6283.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6284 (.I0(\XII[11][4] ), .I1(\XII[9][4] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6284.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6285 (.I0(\XII[10][4] ), .I1(\XII[8][4] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6285.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6286 (.I0(\INSTRUCTION[17] ), .I1(n4648), .I2(n4647), 
            .I3(\INSTRUCTION[18] ), .O(n4649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6286.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6287 (.I0(n4646), .I1(n4645), .I2(\INSTRUCTION[17] ), 
            .I3(n4649), .O(n4650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6287.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6288 (.I0(n4644), .I1(\INSTRUCTION[19] ), .I2(n4650), 
            .O(n4651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6288.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6289 (.I0(n3155), .I1(n51750), .I2(n3174), .O(n4652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6289.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6290 (.I0(n4651), .I1(n3155), .I2(n4639), .I3(n4652), 
            .O(n570_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6290.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6291 (.I0(\XII[26][3] ), .I1(\XII[24][3] ), .I2(\INSTRUCTION[16] ), 
            .O(n4653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6291.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6292 (.I0(\XII[18][3] ), .I1(\XII[16][3] ), .I2(\INSTRUCTION[16] ), 
            .O(n4654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6292.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6293 (.I0(n4654), .I1(n4653), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[18] ), .O(n4655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6293.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6294 (.I0(\XII[17][3] ), .I1(\XII[19][3] ), .I2(n51786), 
            .O(n4656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6294.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6295 (.I0(\XII[25][3] ), .I1(\XII[27][3] ), .I2(n51786), 
            .O(n4657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6295.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6296 (.I0(n4657), .I1(n4656), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6296.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6297 (.I0(\XII[22][3] ), .I1(\XII[20][3] ), .I2(\INSTRUCTION[16] ), 
            .O(n4659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6297.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6298 (.I0(\XII[23][3] ), .I1(\XII[21][3] ), .I2(\INSTRUCTION[16] ), 
            .O(n4660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6298.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6299 (.I0(n4660), .I1(n4659), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6299.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6300 (.I0(\XII[30][3] ), .I1(\XII[28][3] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6300.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6301 (.I0(\XII[31][3] ), .I1(\XII[29][3] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6301.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6302 (.I0(n4662), .I1(n4663), .I2(\INSTRUCTION[18] ), 
            .O(n4664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6302.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6303 (.I0(n4664), .I1(n4661), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[19] ), .O(n4665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6303.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6304 (.I0(n4658), .I1(\INSTRUCTION[17] ), .I2(n4655), 
            .I3(n4665), .O(n4666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6304.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6305 (.I0(\XII[3][3] ), .I1(\XII[1][3] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6305.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6306 (.I0(\XII[2][3] ), .I1(\XII[0][3] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4667), .O(n4668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6306.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6307 (.I0(\XII[7][3] ), .I1(\XII[5][3] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6307.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6308 (.I0(\XII[6][3] ), .I1(\XII[4][3] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4669), .O(n4670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6308.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6309 (.I0(n4670), .I1(n4668), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6309.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6310 (.I0(\XII[15][3] ), .I1(\XII[13][3] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6310.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6311 (.I0(\XII[14][3] ), .I1(\XII[12][3] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6311.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6312 (.I0(\XII[11][3] ), .I1(\XII[9][3] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6312.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6313 (.I0(\XII[10][3] ), .I1(\XII[8][3] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6313.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6314 (.I0(\INSTRUCTION[17] ), .I1(n4675), .I2(n4674), 
            .I3(\INSTRUCTION[18] ), .O(n4676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6314.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6315 (.I0(n4673), .I1(n4672), .I2(\INSTRUCTION[17] ), 
            .I3(n4676), .O(n4677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6315.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6316 (.I0(n4671), .I1(\INSTRUCTION[19] ), .I2(n4677), 
            .O(n4678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6316.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6317 (.I0(n3155), .I1(n51754), .I2(n3174), .O(n4679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6317.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6318 (.I0(n4678), .I1(n3155), .I2(n4666), .I3(n4679), 
            .O(n571_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6318.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6319 (.I0(\XII[26][2] ), .I1(\XII[24][2] ), .I2(\INSTRUCTION[16] ), 
            .O(n4680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6319.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6320 (.I0(\XII[18][2] ), .I1(\XII[16][2] ), .I2(\INSTRUCTION[16] ), 
            .O(n4681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6320.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6321 (.I0(n4681), .I1(n4680), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[18] ), .O(n4682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6321.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6322 (.I0(\XII[17][2] ), .I1(\XII[19][2] ), .I2(n51786), 
            .O(n4683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6322.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6323 (.I0(\XII[25][2] ), .I1(\XII[27][2] ), .I2(n51786), 
            .O(n4684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6323.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6324 (.I0(n4684), .I1(n4683), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6324.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6325 (.I0(\XII[22][2] ), .I1(\XII[20][2] ), .I2(\INSTRUCTION[16] ), 
            .O(n4686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6325.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6326 (.I0(\XII[23][2] ), .I1(\XII[21][2] ), .I2(\INSTRUCTION[16] ), 
            .O(n4687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6326.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6327 (.I0(n4687), .I1(n4686), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6327.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6328 (.I0(\XII[30][2] ), .I1(\XII[28][2] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6328.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6329 (.I0(\XII[31][2] ), .I1(\XII[29][2] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6329.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6330 (.I0(n4689), .I1(n4690), .I2(\INSTRUCTION[18] ), 
            .O(n4691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6330.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6331 (.I0(n4691), .I1(n4688), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[19] ), .O(n4692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6331.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6332 (.I0(n4685), .I1(\INSTRUCTION[17] ), .I2(n4682), 
            .I3(n4692), .O(n4693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6332.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6333 (.I0(\XII[3][2] ), .I1(\XII[1][2] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6333.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6334 (.I0(\XII[2][2] ), .I1(\XII[0][2] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4694), .O(n4695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6334.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6335 (.I0(\XII[7][2] ), .I1(\XII[5][2] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6335.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6336 (.I0(\XII[6][2] ), .I1(\XII[4][2] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4696), .O(n4697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6336.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6337 (.I0(n4697), .I1(n4695), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6337.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6338 (.I0(\XII[15][2] ), .I1(\XII[13][2] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6338.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6339 (.I0(\XII[14][2] ), .I1(\XII[12][2] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6339.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6340 (.I0(\XII[11][2] ), .I1(\XII[9][2] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6340.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6341 (.I0(\XII[10][2] ), .I1(\XII[8][2] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6341.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6342 (.I0(\INSTRUCTION[17] ), .I1(n4702), .I2(n4701), 
            .I3(\INSTRUCTION[18] ), .O(n4703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6342.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6343 (.I0(n4700), .I1(n4699), .I2(\INSTRUCTION[17] ), 
            .I3(n4703), .O(n4704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6343.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6344 (.I0(n4698), .I1(\INSTRUCTION[19] ), .I2(n4704), 
            .O(n4705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6344.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6345 (.I0(n3155), .I1(n51758), .I2(n3174), .O(n4706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6345.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6346 (.I0(n4705), .I1(n3155), .I2(n4693), .I3(n4706), 
            .O(n572_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6346.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6347 (.I0(\XII[3][1] ), .I1(\XII[1][1] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6347.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6348 (.I0(\XII[0][1] ), .I1(\XII[2][1] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4707), .O(n4708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__6348.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__6349 (.I0(\XII[7][1] ), .I1(\XII[5][1] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6349.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6350 (.I0(\XII[6][1] ), .I1(\XII[4][1] ), .I2(\INSTRUCTION[15] ), 
            .I3(n4709), .O(n4710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6350.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6351 (.I0(n4710), .I1(n4708), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[17] ), .O(n4711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__6351.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__6352 (.I0(\XII[15][1] ), .I1(\XII[13][1] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6352.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6353 (.I0(\XII[14][1] ), .I1(\XII[12][1] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6353.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6354 (.I0(\XII[11][1] ), .I1(\XII[9][1] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6354.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6355 (.I0(\XII[10][1] ), .I1(\XII[8][1] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6355.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6356 (.I0(\INSTRUCTION[17] ), .I1(n4715), .I2(n4714), 
            .I3(\INSTRUCTION[18] ), .O(n4716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6356.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6357 (.I0(n4713), .I1(n4712), .I2(\INSTRUCTION[17] ), 
            .I3(n4716), .O(n4717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6357.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6358 (.I0(\INSTRUCTION[19] ), .I1(n4711), .I2(n4717), 
            .I3(n3155), .O(n4718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__6358.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__6359 (.I0(\XII[18][1] ), .I1(\XII[16][1] ), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[16] ), .O(n4719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6359.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6360 (.I0(\XII[26][1] ), .I1(\XII[24][1] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[18] ), .O(n4720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6360.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6361 (.I0(\XII[27][1] ), .I1(\XII[19][1] ), .I2(n51786), 
            .I3(\INSTRUCTION[18] ), .O(n4721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6361.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6362 (.I0(\XII[25][1] ), .I1(\XII[17][1] ), .I2(n51786), 
            .I3(n4721), .O(n4722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6362.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6363 (.I0(n4720), .I1(n4719), .I2(n4722), .I3(\INSTRUCTION[15] ), 
            .O(n4723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6363.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6364 (.I0(\XII[30][1] ), .I1(\XII[28][1] ), .I2(\INSTRUCTION[15] ), 
            .I3(\INSTRUCTION[16] ), .O(n4724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6364.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6365 (.I0(\XII[31][1] ), .I1(\XII[29][1] ), .I2(\INSTRUCTION[16] ), 
            .I3(\INSTRUCTION[15] ), .O(n4725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6365.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6366 (.I0(\XII[22][1] ), .I1(\XII[20][1] ), .I2(\INSTRUCTION[16] ), 
            .O(n4726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6366.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6367 (.I0(\XII[23][1] ), .I1(\XII[21][1] ), .I2(\INSTRUCTION[16] ), 
            .O(n4727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6367.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6368 (.I0(n4727), .I1(n4726), .I2(\INSTRUCTION[18] ), 
            .I3(\INSTRUCTION[15] ), .O(n4728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6368.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6369 (.I0(n4725), .I1(n4724), .I2(\INSTRUCTION[18] ), 
            .I3(n4728), .O(n4729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6369.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6370 (.I0(n4729), .I1(n4723), .I2(\INSTRUCTION[17] ), 
            .I3(\INSTRUCTION[19] ), .O(n4730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6370.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6371 (.I0(n3155), .I1(n51762), .I2(n3174), .O(n4731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6371.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6372 (.I0(n4730), .I1(n4718), .I2(n4731), .O(n573_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6372.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6373 (.I0(n1615_2), .I1(\LOAD_DATA[0] ), .I2(LOAD_OP), 
            .O(n19664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6373.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6374 (.I0(\GPR[0] ), .I1(\GPR[1] ), .O(n4732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6374.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6375 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(\GPR[4] ), .I3(n4732), 
            .O(n4733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6375.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6376 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4733), .O(ceg_net27233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6376.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6377 (.I0(\GPR[1] ), .I1(\GPR[0] ), .O(n4734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6377.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6378 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(\GPR[4] ), .I3(n4734), 
            .O(n4735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6378.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6379 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4735), .O(ceg_net27485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6379.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6380 (.I0(\GPR[0] ), .I1(\GPR[1] ), .O(n4736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6380.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6381 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(\GPR[4] ), .I3(n4736), 
            .O(n4737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6381.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6382 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4737), .O(ceg_net27737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6382.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6383 (.I0(\GPR[0] ), .I1(\GPR[1] ), .O(n4738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6383.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6384 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(\GPR[4] ), .I3(n4738), 
            .O(n4739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6384.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6385 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4739), .O(ceg_net27989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6385.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6386 (.I0(\GPR[3] ), .I1(\GPR[4] ), .I2(n4732), .I3(\GPR[2] ), 
            .O(n4740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6386.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6387 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4740), .O(ceg_net28241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6387.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6388 (.I0(\GPR[3] ), .I1(\GPR[4] ), .I2(n4734), .I3(\GPR[2] ), 
            .O(n4741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6388.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6389 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4741), .O(ceg_net28493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6389.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6390 (.I0(\GPR[3] ), .I1(\GPR[4] ), .I2(n4736), .I3(\GPR[2] ), 
            .O(n4742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6390.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6391 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4742), .O(ceg_net28745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6391.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6392 (.I0(\GPR[3] ), .I1(\GPR[4] ), .I2(n4738), .I3(\GPR[2] ), 
            .O(n4743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6392.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6393 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4743), .O(ceg_net28997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6393.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6394 (.I0(\GPR[2] ), .I1(\GPR[4] ), .I2(\GPR[3] ), .I3(n4732), 
            .O(n4744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6394.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6395 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4744), .O(ceg_net29249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6395.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6396 (.I0(\GPR[2] ), .I1(\GPR[4] ), .I2(\GPR[3] ), .I3(n4734), 
            .O(n4745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6396.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6397 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4745), .O(ceg_net29501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6397.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6398 (.I0(\GPR[2] ), .I1(\GPR[4] ), .I2(\GPR[3] ), .I3(n4736), 
            .O(n4746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6398.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6399 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4746), .O(ceg_net29753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6399.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6400 (.I0(\GPR[2] ), .I1(\GPR[4] ), .I2(\GPR[3] ), .I3(n4738), 
            .O(n4747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6400.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6401 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4747), .O(ceg_net30005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6401.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6402 (.I0(\GPR[4] ), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(n4732), 
            .O(n4748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6402.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6403 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4748), .O(ceg_net30257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6403.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6404 (.I0(\GPR[4] ), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(n4734), 
            .O(n4749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6404.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6405 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4749), .O(ceg_net30509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6405.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6406 (.I0(\GPR[4] ), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(n4736), 
            .O(n4750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6406.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6407 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4750), .O(ceg_net30761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6407.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6408 (.I0(\GPR[4] ), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(n4738), 
            .O(n4751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6408.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6409 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4751), .O(ceg_net31013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6409.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6410 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(n4732), .I3(\GPR[4] ), 
            .O(n4752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6410.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6411 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4752), .O(ceg_net31265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6411.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6412 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(n4734), .I3(\GPR[4] ), 
            .O(n4753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6412.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6413 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4753), .O(ceg_net31517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6413.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6414 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(n4736), .I3(\GPR[4] ), 
            .O(n4754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6414.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6415 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4754), .O(ceg_net31769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6415.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6416 (.I0(\GPR[2] ), .I1(\GPR[3] ), .I2(n4738), .I3(\GPR[4] ), 
            .O(n4755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6416.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6417 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4755), .O(ceg_net32021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6417.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6418 (.I0(\GPR[3] ), .I1(\GPR[2] ), .I2(n4732), .I3(\GPR[4] ), 
            .O(n4756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6418.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6419 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4756), .O(ceg_net32273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6419.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6420 (.I0(\GPR[3] ), .I1(\GPR[2] ), .I2(n4734), .I3(\GPR[4] ), 
            .O(n4757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6420.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6421 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4757), .O(ceg_net32525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6421.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6422 (.I0(\GPR[3] ), .I1(\GPR[2] ), .I2(n4736), .I3(\GPR[4] ), 
            .O(n4758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6422.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6423 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4758), .O(ceg_net32777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6423.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6424 (.I0(\GPR[3] ), .I1(\GPR[2] ), .I2(n4738), .I3(\GPR[4] ), 
            .O(n4759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6424.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6425 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4759), .O(ceg_net33029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6425.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6426 (.I0(\GPR[2] ), .I1(n4732), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6426.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6427 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4760), .O(ceg_net33281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6427.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6428 (.I0(\GPR[2] ), .I1(n4734), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6428.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6429 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4761), .O(ceg_net33533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6429.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6430 (.I0(\GPR[2] ), .I1(n4736), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6430.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6431 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4762), .O(ceg_net33785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6431.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6432 (.I0(\GPR[2] ), .I1(n4738), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6432.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6433 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4763), .O(ceg_net34037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6433.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6434 (.I0(n4732), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6434.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6435 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4764), .O(ceg_net34289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6435.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6436 (.I0(n4734), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6436.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6437 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4765), .O(ceg_net34541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6437.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6438 (.I0(n4736), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6438.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6439 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4766), .O(ceg_net34793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6439.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6440 (.I0(n4738), .I1(\GPR[2] ), .I2(\GPR[3] ), .I3(\GPR[4] ), 
            .O(n4767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6440.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6441 (.I0(MEM_STORE), .I1(STAGE4_EN), .I2(n4767), .O(ceg_net18979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6441.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6442 (.I0(\XI[7][20] ), .I1(\XI[6][20] ), .I2(n2954), 
            .I3(n2953), .O(n4768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6442.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6443 (.I0(\XI[5][20] ), .I1(\XI[4][20] ), .I2(n2953), 
            .I3(n2954), .O(n4769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6443.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6444 (.I0(\XI[3][20] ), .I1(\XI[1][20] ), .I2(n2954), 
            .I3(n2953), .O(n4770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6444.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6445 (.I0(\XI[2][20] ), .I1(\XI[0][20] ), .I2(n2954), 
            .I3(n4770), .O(n4771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6445.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6446 (.I0(n4769), .I1(n4768), .I2(n4771), .I3(n2959), 
            .O(n4772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6446.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6447 (.I0(\XI[15][20] ), .I1(\XI[14][20] ), .I2(n2954), 
            .I3(n2953), .O(n4773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6447.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6448 (.I0(\XI[13][20] ), .I1(\XI[12][20] ), .I2(n2953), 
            .I3(n2954), .O(n4774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6448.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6449 (.I0(\XI[11][20] ), .I1(\XI[9][20] ), .I2(n2954), 
            .I3(n2953), .O(n4775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6449.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6450 (.I0(\XI[10][20] ), .I1(\XI[8][20] ), .I2(n2954), 
            .I3(n4775), .O(n4776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6450.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6451 (.I0(n4774), .I1(n4773), .I2(n4776), .I3(n2959), 
            .O(n4777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6451.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6452 (.I0(n4777), .I1(n4772), .I2(n2966), .I3(n2967), 
            .O(n4778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6452.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6453 (.I0(\XI[19][20] ), .I1(\XI[17][20] ), .I2(n2954), 
            .I3(n2953), .O(n4779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6453.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6454 (.I0(\XI[18][20] ), .I1(\XI[16][20] ), .I2(n2954), 
            .I3(n4779), .O(n4780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6454.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6455 (.I0(\XI[23][20] ), .I1(\XI[21][20] ), .I2(n2954), 
            .I3(n2953), .O(n4781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6455.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6456 (.I0(\XI[22][20] ), .I1(\XI[20][20] ), .I2(n2954), 
            .I3(n4781), .O(n4782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6456.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6457 (.I0(n4782), .I1(n4780), .I2(n2967), .I3(n2959), 
            .O(n4783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6457.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6458 (.I0(\XI[27][20] ), .I1(\XI[26][20] ), .I2(n2954), 
            .I3(n2953), .O(n4784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6458.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6459 (.I0(\XI[25][20] ), .I1(\XI[24][20] ), .I2(n2953), 
            .I3(n2954), .O(n4785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6459.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6460 (.I0(\XI[31][20] ), .I1(\XI[30][20] ), .I2(n2954), 
            .I3(n2953), .O(n4786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6460.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6461 (.I0(\XI[29][20] ), .I1(\XI[28][20] ), .I2(n2953), 
            .I3(n2954), .O(n4787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6461.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6462 (.I0(n4787), .I1(n4786), .I2(n2959), .I3(n2967), 
            .O(n4788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6462.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6463 (.I0(n4785), .I1(n2959), .I2(n4784), .I3(n4788), 
            .O(n4789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6463.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6464 (.I0(n4783), .I1(n4789), .I2(n2966), .O(n4790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6464.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6465 (.I0(n2983), .I1(\PC[20] ), .I2(n2986), .O(n4791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6465.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6466 (.I0(\PC[20] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n4792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6466.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6467 (.I0(n4792), .I1(n3029), .I2(n4791), .I3(n2991), 
            .O(n4793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6467.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6468 (.I0(n4790), .I1(n4778), .I2(n2987), .I3(n4793), 
            .O(n506_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__6468.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__6469 (.I0(\XI[7][29] ), .I1(\XI[6][29] ), .I2(n2954), 
            .I3(n2953), .O(n4794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6469.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6470 (.I0(\XI[5][29] ), .I1(\XI[4][29] ), .I2(n2953), 
            .I3(n2954), .O(n4795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6470.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6471 (.I0(\XI[3][29] ), .I1(\XI[1][29] ), .I2(n2954), 
            .I3(n2953), .O(n4796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6471.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6472 (.I0(\XI[2][29] ), .I1(\XI[0][29] ), .I2(n2954), 
            .I3(n4796), .O(n4797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6472.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6473 (.I0(n4795), .I1(n4794), .I2(n4797), .I3(n2959), 
            .O(n4798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6473.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6474 (.I0(\XI[15][29] ), .I1(\XI[14][29] ), .I2(n2954), 
            .I3(n2953), .O(n4799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6474.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6475 (.I0(\XI[13][29] ), .I1(\XI[12][29] ), .I2(n2953), 
            .I3(n2954), .O(n4800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6475.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6476 (.I0(\XI[11][29] ), .I1(\XI[9][29] ), .I2(n2954), 
            .I3(n2953), .O(n4801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6476.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6477 (.I0(\XI[10][29] ), .I1(\XI[8][29] ), .I2(n2954), 
            .I3(n4801), .O(n4802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6477.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6478 (.I0(n4800), .I1(n4799), .I2(n4802), .I3(n2959), 
            .O(n4803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6478.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6479 (.I0(n4803), .I1(n4798), .I2(n2966), .I3(n2967), 
            .O(n4804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6479.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6480 (.I0(\XI[19][29] ), .I1(\XI[17][29] ), .I2(n2954), 
            .I3(n2953), .O(n4805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6480.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6481 (.I0(\XI[18][29] ), .I1(\XI[16][29] ), .I2(n2954), 
            .I3(n4805), .O(n4806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6481.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6482 (.I0(\XI[23][29] ), .I1(\XI[21][29] ), .I2(n2954), 
            .I3(n2953), .O(n4807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6482.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6483 (.I0(\XI[22][29] ), .I1(\XI[20][29] ), .I2(n2954), 
            .I3(n4807), .O(n4808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6483.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6484 (.I0(n4808), .I1(n4806), .I2(n2967), .I3(n2959), 
            .O(n4809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6484.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6485 (.I0(\XI[27][29] ), .I1(\XI[26][29] ), .I2(n2954), 
            .I3(n2953), .O(n4810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6485.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6486 (.I0(\XI[25][29] ), .I1(\XI[24][29] ), .I2(n2953), 
            .I3(n2954), .O(n4811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6486.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6487 (.I0(\XI[31][29] ), .I1(\XI[30][29] ), .I2(n2954), 
            .I3(n2953), .O(n4812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6487.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6488 (.I0(\XI[29][29] ), .I1(\XI[28][29] ), .I2(n2953), 
            .I3(n2954), .O(n4813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6488.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6489 (.I0(n4813), .I1(n4812), .I2(n2959), .I3(n2967), 
            .O(n4814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6489.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6490 (.I0(n4811), .I1(n2959), .I2(n4810), .I3(n4814), 
            .O(n4815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6490.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6491 (.I0(n4809), .I1(n4815), .I2(n2966), .O(n4816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6491.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6492 (.I0(n2983), .I1(\PC[29] ), .I2(n2986), .O(n4817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6492.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6493 (.I0(\PC[29] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n4818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6493.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6494 (.I0(n4818), .I1(n3029), .I2(n4817), .I3(n2991), 
            .O(n4819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6494.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6495 (.I0(n4816), .I1(n4804), .I2(n2987), .I3(n4819), 
            .O(n497_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__6495.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__6496 (.I0(\XI[7][28] ), .I1(\XI[6][28] ), .I2(n2954), 
            .I3(n2953), .O(n4820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6496.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6497 (.I0(\XI[5][28] ), .I1(\XI[4][28] ), .I2(n2953), 
            .I3(n2954), .O(n4821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6497.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6498 (.I0(\XI[3][28] ), .I1(\XI[1][28] ), .I2(n2954), 
            .I3(n2953), .O(n4822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6498.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6499 (.I0(\XI[2][28] ), .I1(\XI[0][28] ), .I2(n2954), 
            .I3(n4822), .O(n4823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6499.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6500 (.I0(n4821), .I1(n4820), .I2(n4823), .I3(n2959), 
            .O(n4824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6500.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6501 (.I0(\XI[15][28] ), .I1(\XI[14][28] ), .I2(n2954), 
            .I3(n2953), .O(n4825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6501.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6502 (.I0(\XI[13][28] ), .I1(\XI[12][28] ), .I2(n2953), 
            .I3(n2954), .O(n4826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6502.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6503 (.I0(\XI[11][28] ), .I1(\XI[9][28] ), .I2(n2954), 
            .I3(n2953), .O(n4827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6503.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6504 (.I0(\XI[10][28] ), .I1(\XI[8][28] ), .I2(n2954), 
            .I3(n4827), .O(n4828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6504.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6505 (.I0(n4826), .I1(n4825), .I2(n4828), .I3(n2959), 
            .O(n4829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6505.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6506 (.I0(n4829), .I1(n4824), .I2(n2966), .I3(n2967), 
            .O(n4830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6506.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6507 (.I0(\XI[19][28] ), .I1(\XI[17][28] ), .I2(n2954), 
            .I3(n2953), .O(n4831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6507.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6508 (.I0(\XI[18][28] ), .I1(\XI[16][28] ), .I2(n2954), 
            .I3(n4831), .O(n4832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6508.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6509 (.I0(\XI[23][28] ), .I1(\XI[21][28] ), .I2(n2954), 
            .I3(n2953), .O(n4833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6509.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6510 (.I0(\XI[22][28] ), .I1(\XI[20][28] ), .I2(n2954), 
            .I3(n4833), .O(n4834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6510.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6511 (.I0(n4834), .I1(n4832), .I2(n2967), .I3(n2959), 
            .O(n4835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6511.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6512 (.I0(\XI[27][28] ), .I1(\XI[26][28] ), .I2(n2954), 
            .I3(n2953), .O(n4836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6512.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6513 (.I0(\XI[25][28] ), .I1(\XI[24][28] ), .I2(n2953), 
            .I3(n2954), .O(n4837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6513.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6514 (.I0(\XI[31][28] ), .I1(\XI[30][28] ), .I2(n2954), 
            .I3(n2953), .O(n4838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6514.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6515 (.I0(\XI[29][28] ), .I1(\XI[28][28] ), .I2(n2953), 
            .I3(n2954), .O(n4839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6515.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6516 (.I0(n4839), .I1(n4838), .I2(n2959), .I3(n2967), 
            .O(n4840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6516.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6517 (.I0(n4837), .I1(n2959), .I2(n4836), .I3(n4840), 
            .O(n4841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6517.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6518 (.I0(n4835), .I1(n4841), .I2(n2966), .O(n4842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6518.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6519 (.I0(n2983), .I1(\PC[28] ), .I2(n2986), .O(n4843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6519.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6520 (.I0(\PC[28] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n4844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6520.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6521 (.I0(n4844), .I1(n3029), .I2(n4843), .I3(n2991), 
            .O(n4845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6521.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6522 (.I0(n4842), .I1(n4830), .I2(n2987), .I3(n4845), 
            .O(n498_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__6522.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__6523 (.I0(\XI[7][27] ), .I1(\XI[6][27] ), .I2(n2954), 
            .I3(n2953), .O(n4846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6523.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6524 (.I0(\XI[5][27] ), .I1(\XI[4][27] ), .I2(n2953), 
            .I3(n2954), .O(n4847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6524.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6525 (.I0(\XI[3][27] ), .I1(\XI[1][27] ), .I2(n2954), 
            .I3(n2953), .O(n4848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6525.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6526 (.I0(\XI[2][27] ), .I1(\XI[0][27] ), .I2(n2954), 
            .I3(n4848), .O(n4849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6526.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6527 (.I0(n4847), .I1(n4846), .I2(n4849), .I3(n2959), 
            .O(n4850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6527.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6528 (.I0(\XI[15][27] ), .I1(\XI[14][27] ), .I2(n2954), 
            .I3(n2953), .O(n4851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6528.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6529 (.I0(\XI[13][27] ), .I1(\XI[12][27] ), .I2(n2953), 
            .I3(n2954), .O(n4852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6529.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6530 (.I0(\XI[11][27] ), .I1(\XI[9][27] ), .I2(n2954), 
            .I3(n2953), .O(n4853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6530.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6531 (.I0(\XI[10][27] ), .I1(\XI[8][27] ), .I2(n2954), 
            .I3(n4853), .O(n4854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6531.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6532 (.I0(n4852), .I1(n4851), .I2(n4854), .I3(n2959), 
            .O(n4855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6532.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6533 (.I0(n4855), .I1(n4850), .I2(n2966), .I3(n2967), 
            .O(n4856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6533.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6534 (.I0(\XI[19][27] ), .I1(\XI[17][27] ), .I2(n2954), 
            .I3(n2953), .O(n4857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6534.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6535 (.I0(\XI[18][27] ), .I1(\XI[16][27] ), .I2(n2954), 
            .I3(n4857), .O(n4858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6535.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6536 (.I0(\XI[23][27] ), .I1(\XI[21][27] ), .I2(n2954), 
            .I3(n2953), .O(n4859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6536.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6537 (.I0(\XI[22][27] ), .I1(\XI[20][27] ), .I2(n2954), 
            .I3(n4859), .O(n4860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6537.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6538 (.I0(n4860), .I1(n4858), .I2(n2967), .I3(n2959), 
            .O(n4861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6538.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6539 (.I0(\XI[27][27] ), .I1(\XI[26][27] ), .I2(n2954), 
            .I3(n2953), .O(n4862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6539.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6540 (.I0(\XI[25][27] ), .I1(\XI[24][27] ), .I2(n2953), 
            .I3(n2954), .O(n4863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6540.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6541 (.I0(\XI[31][27] ), .I1(\XI[30][27] ), .I2(n2954), 
            .I3(n2953), .O(n4864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6541.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6542 (.I0(\XI[29][27] ), .I1(\XI[28][27] ), .I2(n2953), 
            .I3(n2954), .O(n4865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6542.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6543 (.I0(n4865), .I1(n4864), .I2(n2959), .I3(n2967), 
            .O(n4866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6543.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6544 (.I0(n4863), .I1(n2959), .I2(n4862), .I3(n4866), 
            .O(n4867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6544.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6545 (.I0(n4861), .I1(n4867), .I2(n2966), .O(n4868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6545.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6546 (.I0(n2983), .I1(\PC[27] ), .I2(n2986), .O(n4869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6546.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6547 (.I0(\PC[27] ), .I1(n3026), .I2(n3379), .I3(n2986), 
            .O(n4870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6547.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6548 (.I0(n4870), .I1(n3029), .I2(n4869), .I3(n2991), 
            .O(n4871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6548.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6549 (.I0(n4868), .I1(n4856), .I2(n2987), .I3(n4871), 
            .O(n499_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__6549.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__6550 (.I0(n3509), .I1(n3508), .I2(\SHIFT_STEPS[0] ), 
            .O(n4872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6550.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6551 (.I0(\ARG1[4] ), .I1(\ARG1[2] ), .I2(\SHIFT_STEPS[1] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6551.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6552 (.I0(\ARG1[8] ), .I1(\ARG1[6] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6552.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6553 (.I0(n3505), .I1(n4874), .I2(\SHIFT_STEPS[0] ), 
            .O(n4875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6553.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6554 (.I0(n4873), .I1(n4872), .I2(n4875), .I3(\SHIFT_STEPS[2] ), 
            .O(n4876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6554.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6555 (.I0(\ARG1[20] ), .I1(\ARG1[18] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6555.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6556 (.I0(n3531), .I1(n4877), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6556.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6557 (.I0(\ARG1[24] ), .I1(\ARG1[22] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6557.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6558 (.I0(n3528), .I1(n4879), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6558.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6559 (.I0(n4878), .I1(n4880), .O(n4881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6559.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6560 (.I0(n4881), .I1(n4876), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[4] ), .O(n4882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__6560.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__6561 (.I0(\ARG1[28] ), .I1(\ARG1[26] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6561.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6562 (.I0(n3524), .I1(n4883), .I2(\SHIFT_STEPS[0] ), 
            .O(n4884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6562.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6563 (.I0(\ARG1[30] ), .I1(\ARG1[29] ), .I2(\SHIFT_STEPS[0] ), 
            .O(n4885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6563.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6564 (.I0(n4885), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6564.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6565 (.I0(n4886), .I1(n4884), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[4] ), .O(n4887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6565.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6566 (.I0(\ARG1[16] ), .I1(\ARG1[14] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6566.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6567 (.I0(n3513), .I1(n4888), .I2(\SHIFT_STEPS[0] ), 
            .O(n4889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6567.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6568 (.I0(\ARG1[12] ), .I1(\ARG1[10] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6568.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6569 (.I0(n3516), .I1(n4890), .I2(\SHIFT_STEPS[0] ), 
            .O(n4891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6569.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6570 (.I0(n4891), .I1(n4889), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6570.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6571 (.I0(n4892), .I1(n4887), .I2(\SHIFT_STEPS[3] ), 
            .O(n4893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6571.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6572 (.I0(\OPERATION[0] ), .I1(\ARG2[1] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[1] ), .O(n4894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6572.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6573 (.I0(n4894), .I1(\OPERATION[2] ), .O(n4895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6573.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6574 (.I0(n4893), .I1(n4882), .I2(n3536), .I3(n4895), 
            .O(n4896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6574.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6575 (.I0(\ARG1[0] ), .I1(\ARG1[1] ), .I2(\SHIFT_STEPS[1] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6575.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6576 (.I0(n1371), .I1(n1448), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n4898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6576.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6577 (.I0(n3543), .I1(n4897), .I2(n4898), .I3(\OPERATION[2] ), 
            .O(n4899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6577.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6578 (.I0(n4893), .I1(n4882), .I2(n3547), .I3(n4899), 
            .O(n4900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6578.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6579 (.I0(n4896), .I1(n4900), .I2(\OPERATION[3] ), .O(n1614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6579.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6580 (.I0(\ARG1[0] ), .I1(\ARG1[2] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6580.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6581 (.I0(n3508), .I1(n4901), .I2(\SHIFT_STEPS[0] ), 
            .O(n4902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6581.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6582 (.I0(\SHIFT_STEPS[4] ), .I1(n3542), .O(n4903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6582.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6583 (.I0(n4903), .I1(n4902), .I2(n3445), .O(n4904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__6583.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__6584 (.I0(\ARG1[5] ), .I1(\ARG1[3] ), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[1] ), .O(n4905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6584.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6585 (.I0(\ARG1[2] ), .I1(\ARG1[4] ), .I2(\SHIFT_STEPS[0] ), 
            .I3(n4905), .O(n4906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__6585.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__6586 (.I0(\ARG1[9] ), .I1(\ARG1[7] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6586.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6587 (.I0(n4874), .I1(n4907), .I2(\SHIFT_STEPS[0] ), 
            .O(n4908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6587.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6588 (.I0(n4908), .I1(n4906), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6588.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6589 (.I0(\ARG1[17] ), .I1(\ARG1[15] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6589.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6590 (.I0(n4888), .I1(n4910), .I2(\SHIFT_STEPS[0] ), 
            .O(n4911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6590.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6591 (.I0(\ARG1[13] ), .I1(\ARG1[11] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6591.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6592 (.I0(n4890), .I1(n4912), .I2(\SHIFT_STEPS[0] ), 
            .O(n4913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6592.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6593 (.I0(n4913), .I1(n4911), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n4914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6593.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6594 (.I0(\ARG1[25] ), .I1(\ARG1[23] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6594.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6595 (.I0(n4879), .I1(n4915), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6595.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6596 (.I0(\ARG1[21] ), .I1(\ARG1[19] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6596.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6597 (.I0(n4877), .I1(n4917), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6597.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6598 (.I0(\ARG1[28] ), .I1(\ARG1[26] ), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[1] ), .O(n4919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6598.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6599 (.I0(\ARG1[29] ), .I1(\ARG1[27] ), .I2(\SHIFT_STEPS[1] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6599.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6600 (.I0(\ARG1[30] ), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[1] ), .O(n4921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__6600.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__6601 (.I0(n4920), .I1(n4919), .I2(n4921), .I3(\SHIFT_STEPS[2] ), 
            .O(n4922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6601.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6602 (.I0(n4918), .I1(n4916), .I2(n4922), .I3(\SHIFT_STEPS[3] ), 
            .O(n4923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6602.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6603 (.I0(n4914), .I1(n4909), .I2(n4923), .I3(\SHIFT_STEPS[4] ), 
            .O(n4924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6603.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6604 (.I0(n1370), .I1(n1446), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n4925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6604.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6605 (.I0(n4924), .I1(n3547), .I2(n4925), .I3(n3545), 
            .O(n4926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6605.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6606 (.I0(\OPERATION[0] ), .I1(\ARG2[2] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[2] ), .O(n4927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6606.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6607 (.I0(n4924), .I1(n3536), .I2(n4927), .I3(n3537), 
            .O(n4928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6607.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6608 (.I0(n4904), .I1(n4926), .I2(n4928), .O(n1613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__6608.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__6609 (.I0(\OPERATION[0] ), .I1(\ARG2[3] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[3] ), .O(n4929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6609.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6610 (.I0(\ARG1[5] ), .I1(\ARG1[3] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6610.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6611 (.I0(n3506), .I1(n4930), .I2(\SHIFT_STEPS[0] ), 
            .O(n4931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6611.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6612 (.I0(n3517), .I1(n4907), .I2(\SHIFT_STEPS[0] ), 
            .O(n4932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6612.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6613 (.I0(n4932), .I1(n4931), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__6613.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__6614 (.I0(n3532), .I1(n4910), .I2(\SHIFT_STEPS[0] ), 
            .O(n4934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6614.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6615 (.I0(n3514), .I1(n4912), .I2(\SHIFT_STEPS[0] ), 
            .O(n4935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6615.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6616 (.I0(n4935), .I1(n4934), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n4936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6616.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6617 (.I0(\ARG1[29] ), .I1(\ARG1[27] ), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[1] ), .O(n4937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6617.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6618 (.I0(\ARG1[30] ), .I1(\ARG1[28] ), .I2(\SHIFT_STEPS[1] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6618.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6619 (.I0(n4937), .I1(n4938), .I2(\ARG1[31] ), .I3(\SHIFT_STEPS[2] ), 
            .O(n4939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6619.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6620 (.I0(n3529), .I1(n4917), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6620.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6621 (.I0(n3525), .I1(n4915), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6621.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6622 (.I0(n4940), .I1(n4941), .I2(n4939), .I3(\SHIFT_STEPS[3] ), 
            .O(n4942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6622.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6623 (.I0(n4936), .I1(n4933), .I2(n4942), .I3(\SHIFT_STEPS[4] ), 
            .O(n4943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6623.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6624 (.I0(n4943), .I1(n3536), .I2(n4929), .I3(\OPERATION[2] ), 
            .O(n4944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6624.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6625 (.I0(\ARG1[1] ), .I1(\ARG1[3] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6625.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6626 (.I0(n4901), .I1(n4945), .I2(\SHIFT_STEPS[0] ), 
            .O(n4946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6626.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6627 (.I0(n1369), .I1(n1444), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n4947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6627.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6628 (.I0(n3543), .I1(n4946), .I2(n4947), .I3(\OPERATION[2] ), 
            .O(n4948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6628.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6629 (.I0(n4943), .I1(n3547), .I2(n4948), .O(n4949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6629.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6630 (.I0(\RES[3]_2~FF_brt_120_q ), .I1(\RES[3]_2~FF_brt_121_q ), 
            .I2(\RES[4]_2~FF_brt_125_q ), .O(n1612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6630.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6631 (.I0(n3518), .I1(n3507), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6631.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6632 (.I0(n3533), .I1(n3515), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n4951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6632.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6633 (.I0(n3525), .I1(n3524), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6633.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6634 (.I0(n3529), .I1(n3528), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6634.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6635 (.I0(n3521), .I1(n3522), .I2(\ARG1[31] ), .I3(\SHIFT_STEPS[2] ), 
            .O(n4954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6635.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6636 (.I0(n4953), .I1(n4952), .I2(n4954), .I3(\SHIFT_STEPS[3] ), 
            .O(n4955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6636.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6637 (.I0(n4951), .I1(n4950), .I2(n4955), .I3(\SHIFT_STEPS[4] ), 
            .O(n4956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6637.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6638 (.I0(\SHIFT_STEPS[4] ), .I1(n3445), .O(n4957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6638.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6639 (.I0(\SHIFT_STEPS[3] ), .I1(n4957), .O(n4958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6639.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6640 (.I0(\ARG1[2] ), .I1(\ARG1[4] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6640.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6641 (.I0(n4945), .I1(n4959), .I2(\SHIFT_STEPS[0] ), 
            .O(n4960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6641.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6642 (.I0(n4960), .I1(n3541), .I2(\SHIFT_STEPS[2] ), 
            .O(n4961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6642.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6643 (.I0(n1368), .I1(n1442), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n4962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6643.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6644 (.I0(n4961), .I1(n4958), .I2(n4962), .I3(\OPERATION[2] ), 
            .O(n4963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6644.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6645 (.I0(n4956), .I1(n3547), .I2(n4963), .O(n4964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6645.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6646 (.I0(\OPERATION[0] ), .I1(\ARG2[4] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[4] ), .O(n4965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6646.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6647 (.I0(n4956), .I1(n3536), .I2(n4965), .I3(\OPERATION[2] ), 
            .O(n4966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6647.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6648 (.I0(\RES[4]_2~FF_brt_123_q ), .I1(\RES[4]_2~FF_brt_124_q ), 
            .I2(\RES[4]_2~FF_brt_125_q ), .O(n1611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6648.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6649 (.I0(\SHIFT_STEPS[3] ), .I1(\SHIFT_STEPS[4] ), .O(n4967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6649.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6650 (.I0(\ARG1[3] ), .I1(\ARG1[5] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6650.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6651 (.I0(n4959), .I1(n4968), .I2(\SHIFT_STEPS[0] ), 
            .O(n4969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6651.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6652 (.I0(n4969), .I1(n4897), .I2(\SHIFT_STEPS[2] ), 
            .O(n4970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6652.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6653 (.I0(n4970), .I1(n4967), .I2(n3445), .O(n4971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6653.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6654 (.I0(n4891), .I1(n4875), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6654.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6655 (.I0(n3531), .I1(n4877), .I2(\SHIFT_STEPS[0] ), 
            .O(n4973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6655.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6656 (.I0(n4889), .I1(n4973), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n4974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6656.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6657 (.I0(n3528), .I1(n4879), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6657.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6658 (.I0(n3524), .I1(n4883), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6658.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6659 (.I0(n4885), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[1] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccc5 */ ;
    defparam LUT__6659.LUTMASK = 16'hccc5;
    EFX_LUT4 LUT__6660 (.I0(n4976), .I1(n4975), .I2(n4977), .I3(\SHIFT_STEPS[3] ), 
            .O(n4978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6660.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6661 (.I0(n4974), .I1(n4972), .I2(n4978), .I3(\SHIFT_STEPS[4] ), 
            .O(n4979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6661.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6662 (.I0(n1367), .I1(n1440), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n4980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6662.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6663 (.I0(n4979), .I1(n3547), .I2(n4980), .I3(n3545), 
            .O(n4981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6663.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6664 (.I0(\OPERATION[0] ), .I1(\ARG2[5] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[5] ), .O(n4982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6664.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6665 (.I0(n4979), .I1(n3536), .I2(n4982), .I3(n3537), 
            .O(n4983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6665.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6666 (.I0(\RES[5]_2~FF_brt_126_q ), .I1(\RES[5]_2~FF_brt_127_q ), 
            .I2(\RES[5]_2~FF_brt_128_q ), .O(n1610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__6666.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__6667 (.I0(n4913), .I1(n4908), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n4984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6667.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6668 (.I0(n4877), .I1(n4917), .I2(\SHIFT_STEPS[0] ), 
            .O(n4985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6668.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6669 (.I0(n4985), .I1(n4911), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n4986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6669.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6670 (.I0(n4919), .I1(n4920), .I2(\SHIFT_STEPS[2] ), 
            .O(n4987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6670.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6671 (.I0(n4879), .I1(n4915), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n4988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6671.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6672 (.I0(n4921), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[2] ), 
            .O(n4989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6672.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6673 (.I0(n4988), .I1(n4987), .I2(n4989), .I3(\SHIFT_STEPS[3] ), 
            .O(n4990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6673.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6674 (.I0(n4986), .I1(n4984), .I2(n4990), .I3(\SHIFT_STEPS[4] ), 
            .O(n4991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6674.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6675 (.I0(\ARG1[4] ), .I1(\ARG1[6] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n4992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6675.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6676 (.I0(n4968), .I1(n4992), .I2(\SHIFT_STEPS[0] ), 
            .O(n4993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6676.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6677 (.I0(n4902), .I1(n4993), .I2(\SHIFT_STEPS[2] ), 
            .O(n4994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__6677.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__6678 (.I0(n4994), .I1(n4967), .I2(n3445), .O(n4995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6678.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6679 (.I0(n1366), .I1(n1438), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n4996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6679.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6680 (.I0(n4995), .I1(n4996), .I2(n3545), .O(n4997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6680.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6681 (.I0(\OPERATION[0] ), .I1(\ARG2[6] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[6] ), .O(n4998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6681.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6682 (.I0(n4991), .I1(n3536), .I2(n4998), .I3(n3537), 
            .O(n4999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6682.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6683 (.I0(\RES[9]_2~FF_brt_1_brt_24_q ), .I1(\RES[6]_2~FF_brt_129_q ), 
            .I2(\RES[6]_2~FF_brt_130_q ), .I3(\RES[6]_2~FF_brt_131_q ), 
            .O(n1609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__6683.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__6684 (.I0(\OPERATION[0] ), .I1(\OPERATION[2] ), .O(n5000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6684.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6685 (.I0(\ARG1[5] ), .I1(\ARG1[7] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6685.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6686 (.I0(n4992), .I1(n5001), .I2(\SHIFT_STEPS[0] ), 
            .O(n5002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6686.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6687 (.I0(n4946), .I1(n5002), .I2(\SHIFT_STEPS[2] ), 
            .O(n5003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6687.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6688 (.I0(n5003), .I1(n4967), .I2(n1436), .I3(\OPERATION[1] ), 
            .O(n5004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__6688.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__6689 (.I0(\SHIFT_STEPS[3] ), .I1(\SHIFT_STEPS[4] ), .O(n5005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6689.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6690 (.I0(n3525), .I1(n4915), .I2(\SHIFT_STEPS[0] ), 
            .O(n5006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6690.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6691 (.I0(n4937), .I1(n4938), .O(n5007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6691.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6692 (.I0(n5007), .I1(n5006), .I2(\SHIFT_STEPS[2] ), 
            .O(n5008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__6692.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__6693 (.I0(\OPERATION[0] ), .I1(\OPERATION[2] ), .I2(\OPERATION[1] ), 
            .O(n5009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6693.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6694 (.I0(n4935), .I1(n4932), .I2(\SHIFT_STEPS[2] ), 
            .I3(n4967), .O(n5010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6694.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6695 (.I0(n5008), .I1(n5005), .I2(n5010), .I3(n5009), 
            .O(n5011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6695.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6696 (.I0(n3529), .I1(n4917), .I2(\SHIFT_STEPS[0] ), 
            .O(n5012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6696.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6697 (.I0(n5012), .I1(n4934), .I2(\SHIFT_STEPS[2] ), 
            .O(n5013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6697.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6698 (.I0(\SHIFT_STEPS[4] ), .I1(\ARG1[31] ), .O(n5014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6698.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6699 (.I0(n5014), .I1(\SHIFT_STEPS[3] ), .O(n5015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6699.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6700 (.I0(n5013), .I1(\SHIFT_STEPS[4] ), .I2(n5015), 
            .O(n5016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6700.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6701 (.I0(\OPERATION[0] ), .I1(\ARG2[7] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[7] ), .O(n5017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6701.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6702 (.I0(\OPERATION[2] ), .I1(\OPERATION[0] ), .O(n5018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6702.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6703 (.I0(\OPERATION[1] ), .I1(n1365), .I2(n5018), .O(n5019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6703.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6704 (.I0(\RES[7]_2~FF_brt_20_brt_70_brt_132_q ), .I1(\RES[17]_2~FF_brt_8_brt_36_q ), 
            .I2(\RES[7]_2~FF_brt_20_brt_70_brt_133_q ), .O(n5020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6704.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6705 (.I0(\RES[7]_2~FF_brt_20_brt_68_q ), .I1(\RES[7]_2~FF_brt_20_brt_69_q ), 
            .I2(n5020), .O(n5021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6705.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6706 (.I0(\RES[7]_2~FF_brt_18_q ), .I1(\RES[7]_2~FF_brt_19_q ), 
            .I2(n5021), .I3(\RES[4]_2~FF_brt_125_q ), .O(n1608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6706.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6707 (.I0(\SHIFT_STEPS[4] ), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[3] ), 
            .O(n5022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__6707.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__6708 (.I0(n3533), .I1(n3530), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n5023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6708.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6709 (.I0(n3518), .I1(n3515), .I2(\SHIFT_STEPS[2] ), 
            .I3(n4967), .O(n5024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6709.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6710 (.I0(n3526), .I1(n3523), .I2(\SHIFT_STEPS[2] ), 
            .I3(n5005), .O(n5025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__6710.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__6711 (.I0(n5023), .I1(n5022), .I2(n5024), .I3(n5025), 
            .O(n5026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6711.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6712 (.I0(\ARG1[6] ), .I1(\ARG1[8] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6712.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6713 (.I0(n5001), .I1(n5027), .I2(\SHIFT_STEPS[0] ), 
            .O(n5028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6713.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6714 (.I0(n4960), .I1(n5028), .I2(\SHIFT_STEPS[2] ), 
            .O(n5029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6714.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6715 (.I0(\SHIFT_STEPS[2] ), .I1(\SHIFT_STEPS[3] ), .O(n5030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6715.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6716 (.I0(n3541), .I1(n5030), .O(n5031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6716.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6717 (.I0(n5029), .I1(\SHIFT_STEPS[3] ), .I2(n5031), 
            .I3(n4957), .O(n5032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__6717.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__6718 (.I0(n1364), .I1(n1434), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n5033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6718.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6719 (.I0(\RES[8]_2~FF_brt_21_brt_73_brt_134_q ), .I1(\RES[17]_2~FF_brt_8_brt_36_q ), 
            .O(n5034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6719.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6720 (.I0(\RES[8]_2~FF_brt_21_brt_71_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(\RES[8]_2~FF_brt_21_brt_72_q ), .I3(n5034), .O(n5035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__6720.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__6721 (.I0(\OPERATION[0] ), .I1(\ARG2[8] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[8] ), .O(n5036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6721.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6722 (.I0(n5026), .I1(n3536), .I2(n5036), .I3(\OPERATION[2] ), 
            .O(n5037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6722.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6723 (.I0(n5035), .I1(\RES[8]_2~FF_brt_22_q ), .I2(\RES[4]_2~FF_brt_125_q ), 
            .O(n1607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6723.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6724 (.I0(n4878), .I1(n4880), .I2(\ARG1[31] ), .I3(\SHIFT_STEPS[4] ), 
            .O(n5038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6724.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6725 (.I0(n4892), .I1(n4887), .I2(n5038), .I3(\SHIFT_STEPS[3] ), 
            .O(n5039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6725.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6726 (.I0(\OPERATION[0] ), .I1(\ARG2[9] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[9] ), .O(n5040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6726.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6727 (.I0(n5039), .I1(n3536), .I2(n5040), .I3(\OPERATION[2] ), 
            .O(n5041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6727.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6728 (.I0(\ARG1[7] ), .I1(\ARG1[9] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6728.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6729 (.I0(n5027), .I1(n5042), .I2(\SHIFT_STEPS[0] ), 
            .O(n5043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6729.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6730 (.I0(n4969), .I1(n5043), .I2(\SHIFT_STEPS[2] ), 
            .O(n5044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6730.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6731 (.I0(n4897), .I1(n5030), .O(n5045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6731.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6732 (.I0(n5044), .I1(\SHIFT_STEPS[3] ), .I2(n5045), 
            .I3(n4957), .O(n5046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__6732.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__6733 (.I0(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_135_q ), 
            .I1(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_q ), .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), 
            .I3(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .O(n5047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6733.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6734 (.I0(n5047), .I1(\RES[17]_2~FF_brt_8_brt_36_q ), 
            .O(n5048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6734.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6735 (.I0(\RES[9]_2~FF_brt_1_brt_23_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(\RES[9]_2~FF_brt_1_brt_25_q ), .I3(n5048), .O(n5049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6735.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6736 (.I0(\RES[9]_2~FF_brt_0_q ), .I1(n5049), .I2(\RES[4]_2~FF_brt_125_q ), 
            .O(n1606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6736.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6737 (.I0(n4918), .I1(n4916), .I2(\SHIFT_STEPS[4] ), 
            .O(n5050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6737.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6738 (.I0(n4922), .I1(n5005), .O(n5051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6738.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6739 (.I0(n4913), .I1(n4911), .I2(\SHIFT_STEPS[2] ), 
            .I3(n4967), .O(n5052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6739.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6740 (.I0(n5050), .I1(n5022), .I2(n5051), .I3(n5052), 
            .O(n5053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6740.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6741 (.I0(\ARG1[8] ), .I1(\ARG1[10] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6741.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6742 (.I0(n5042), .I1(n5054), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[0] ), .O(n5055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6742.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6743 (.I0(n4968), .I1(n4992), .I2(\SHIFT_STEPS[0] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n5056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6743.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6744 (.I0(n3508), .I1(n4901), .I2(\SHIFT_STEPS[0] ), 
            .I3(n5030), .O(n5057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6744.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6745 (.I0(n5056), .I1(\SHIFT_STEPS[3] ), .I2(n5055), 
            .I3(n5057), .O(n5058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__6745.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__6746 (.I0(\RES[10]_2~FF_brt_3_brt_28_brt_76_brt_139_q ), 
            .I1(\RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140_q ), .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), 
            .I3(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .O(n5059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6746.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6747 (.I0(\RES[10]_2~FF_brt_3_brt_28_brt_75_q ), .I1(\RES[17]_2~FF_brt_8_brt_34_q ), 
            .I2(n5059), .I3(\RES[17]_2~FF_brt_8_brt_36_q ), .O(n5060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6747.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6748 (.I0(\RES[10]_2~FF_brt_3_brt_27_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(n5060), .O(n5061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6748.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6749 (.I0(\OPERATION[0] ), .I1(\ARG2[10] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[10] ), .O(n5062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6749.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6750 (.I0(n5053), .I1(n3536), .I2(n5062), .I3(\OPERATION[2] ), 
            .O(n5063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6750.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6751 (.I0(n5061), .I1(\RES[10]_2~FF_brt_4_q ), .I2(\RES[4]_2~FF_brt_125_q ), 
            .O(n1605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6751.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6752 (.I0(\ARG1[9] ), .I1(\ARG1[11] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6752.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6753 (.I0(n5054), .I1(n5064), .I2(\SHIFT_STEPS[0] ), 
            .O(n5065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6753.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6754 (.I0(n5002), .I1(n5065), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n5066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6754.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6755 (.I0(n4946), .I1(n5030), .I2(n5066), .O(n5067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6755.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6756 (.I0(n5067), .I1(n3445), .O(n5068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6756.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6757 (.I0(n4935), .I1(n4934), .I2(\SHIFT_STEPS[2] ), 
            .I3(n4967), .O(n5069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6757.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6758 (.I0(n5007), .I1(\ARG1[31] ), .I2(n3542), .I3(\SHIFT_STEPS[4] ), 
            .O(n5070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6758.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6759 (.I0(\SHIFT_STEPS[4] ), .I1(\SHIFT_STEPS[3] ), .O(n5071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6759.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6760 (.I0(n4940), .I1(n4941), .I2(n5071), .O(n5072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6760.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6761 (.I0(n5069), .I1(n5070), .I2(n5072), .O(n5073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6761.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6762 (.I0(n5073), .I1(n3547), .O(n5074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6762.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6763 (.I0(n3445), .I1(\SHIFT_STEPS[4] ), .O(n5075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6763.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6764 (.I0(n1361), .I1(n1428), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n5076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6764.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6765 (.I0(n5075), .I1(n5076), .I2(n3545), .O(n5077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6765.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6766 (.I0(\OPERATION[0] ), .I1(\ARG2[11] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[11] ), .O(n5078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6766.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6767 (.I0(n5073), .I1(n3536), .I2(n5078), .I3(n3537), 
            .O(n5079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6767.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6768 (.I0(\RES[11]_2~FF_brt_141_q ), .I1(\RES[11]_2~FF_brt_142_q ), 
            .I2(\RES[11]_2~FF_brt_143_q ), .I3(\RES[11]_2~FF_brt_144_q ), 
            .O(n1604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__6768.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__6769 (.I0(\ARG1[10] ), .I1(\ARG1[12] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6769.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6770 (.I0(n5064), .I1(n5080), .I2(\SHIFT_STEPS[0] ), 
            .O(n5081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6770.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6771 (.I0(n5028), .I1(n5081), .I2(\SHIFT_STEPS[2] ), 
            .O(n5082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6771.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6772 (.I0(n4961), .I1(n5082), .I2(\SHIFT_STEPS[3] ), 
            .I3(n3445), .O(n5083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6772.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6773 (.I0(n1360), .I1(n1426), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n5084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6773.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6774 (.I0(\RES[27]_2~FF_brt_53_q ), .I1(\RES[12]_2~FF_brt_78_brt_145_q ), 
            .I2(\RES[4]_2~FF_brt_125_q ), .O(n5085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6774.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6775 (.I0(n5018), .I1(\OPERATION[1] ), .O(n5086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6775.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6776 (.I0(n4953), .I1(n4952), .I2(n5071), .O(n5087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6776.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6777 (.I0(n3523), .I1(\ARG1[31] ), .I2(n3542), .I3(\SHIFT_STEPS[4] ), 
            .O(n5088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6777.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6778 (.I0(n3533), .I1(n3515), .I2(\SHIFT_STEPS[2] ), 
            .I3(n4967), .O(n5089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6778.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6779 (.I0(n5087), .I1(n5088), .I2(n5089), .O(n5090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6779.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6780 (.I0(\OPERATION[0] ), .I1(\ARG2[12] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[12] ), .O(n5091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6780.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6781 (.I0(n5091), .I1(\OPERATION[2] ), .O(n5092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6781.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6782 (.I0(n5086), .I1(n3536), .I2(n5090), .I3(n5092), 
            .O(n5093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c5f */ ;
    defparam LUT__6782.LUTMASK = 16'h0c5f;
    EFX_LUT4 LUT__6783 (.I0(\RES[12]_2~FF_brt_77_q ), .I1(n5085), .I2(\RES[24]_2~FF_brt_48_q ), 
            .I3(\RES[12]_2~FF_brt_79_q ), .O(n1603_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6783.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6784 (.I0(n4975), .I1(\SHIFT_STEPS[4] ), .I2(n4976), 
            .I3(n5015), .O(n5094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6784.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6785 (.I0(n3547), .I1(n3536), .I2(n5094), .I3(\OPERATION[2] ), 
            .O(n5095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6785.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6786 (.I0(n4889), .I1(n4973), .I2(\SHIFT_STEPS[2] ), 
            .O(n5096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6786.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6787 (.I0(n5096), .I1(n4977), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[4] ), .O(n5097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__6787.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__6788 (.I0(\OPERATION[0] ), .I1(\ARG2[13] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[13] ), .O(n5098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6788.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6789 (.I0(n5098), .I1(n5097), .I2(n5095), .I3(\OPERATION[2] ), 
            .O(n5099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h75cf */ ;
    defparam LUT__6789.LUTMASK = 16'h75cf;
    EFX_LUT4 LUT__6790 (.I0(\ARG1[11] ), .I1(\ARG1[13] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6790.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6791 (.I0(n5080), .I1(n5100), .I2(\SHIFT_STEPS[0] ), 
            .O(n5101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6791.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6792 (.I0(n5043), .I1(n5101), .I2(\SHIFT_STEPS[2] ), 
            .O(n5102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6792.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6793 (.I0(n4970), .I1(n5102), .I2(\SHIFT_STEPS[3] ), 
            .O(n5103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6793.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6794 (.I0(n1359), .I1(n1424), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n5104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6794.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6795 (.I0(n5103), .I1(n4957), .I2(n5104), .O(n5105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6795.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6796 (.I0(\RES[13]_2~FF_brt_146_q ), .I1(\RES[17]_2~FF_brt_8_brt_36_q ), 
            .I2(\RES[4]_2~FF_brt_125_q ), .I3(\RES[13]_2~FF_brt_147_q ), 
            .O(n1602_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d03 */ ;
    defparam LUT__6796.LUTMASK = 16'h0d03;
    EFX_LUT4 LUT__6797 (.I0(\ARG1[12] ), .I1(\ARG1[14] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6797.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6798 (.I0(n5100), .I1(n5106), .I2(\SHIFT_STEPS[0] ), 
            .O(n5107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6798.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6799 (.I0(n5042), .I1(n5054), .I2(\SHIFT_STEPS[0] ), 
            .O(n5108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6799.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6800 (.I0(n5108), .I1(n5107), .I2(\SHIFT_STEPS[2] ), 
            .O(n5109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6800.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6801 (.I0(n4994), .I1(n5109), .I2(\SHIFT_STEPS[3] ), 
            .O(n5110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6801.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6802 (.I0(n4985), .I1(n4911), .I2(\SHIFT_STEPS[2] ), 
            .I3(n4967), .O(n5111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6802.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6803 (.I0(n4988), .I1(n4987), .I2(n5071), .O(n5112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6803.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6804 (.I0(n4921), .I1(\ARG1[31] ), .I2(n3542), .I3(\SHIFT_STEPS[4] ), 
            .O(n5113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6804.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6805 (.I0(n5111), .I1(n5112), .I2(n5113), .I3(n3547), 
            .O(n5114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6805.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6806 (.I0(n1358), .I1(n1422), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n5115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6806.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6807 (.I0(n5114), .I1(n5075), .I2(n5115), .I3(n3545), 
            .O(n5116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6807.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6808 (.I0(n5111), .I1(n5112), .I2(n5113), .O(n5117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6808.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6809 (.I0(\OPERATION[0] ), .I1(\ARG2[14] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[14] ), .O(n5118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6809.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6810 (.I0(n5117), .I1(n3536), .I2(n5118), .I3(n3537), 
            .O(n5119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6810.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6811 (.I0(\RES[14]_2~FF_brt_148_q ), .I1(\RES[28]_2~FF_brt_15_brt_59_q ), 
            .I2(\RES[14]_2~FF_brt_149_q ), .I3(\RES[14]_2~FF_brt_150_q ), 
            .O(n1601_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__6811.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__6812 (.I0(n5007), .I1(n5006), .I2(\SHIFT_STEPS[2] ), 
            .I3(n5071), .O(n5120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6812.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6813 (.I0(n5013), .I1(n4967), .I2(n5120), .I3(n5014), 
            .O(n5121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6813.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6814 (.I0(\OPERATION[0] ), .I1(\ARG2[15] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[15] ), .O(n5122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6814.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6815 (.I0(n5121), .I1(n3536), .I2(n5122), .I3(\OPERATION[2] ), 
            .O(n5123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6815.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6816 (.I0(\ARG1[13] ), .I1(\ARG1[15] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6816.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6817 (.I0(n5106), .I1(n5124), .I2(\SHIFT_STEPS[0] ), 
            .O(n5125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6817.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6818 (.I0(n5065), .I1(n5125), .I2(\SHIFT_STEPS[2] ), 
            .O(n5126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6818.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6819 (.I0(n5003), .I1(n5126), .I2(\SHIFT_STEPS[3] ), 
            .I3(n4957), .O(n5127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6819.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6820 (.I0(n1357), .I1(n1420), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n5128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6820.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6821 (.I0(\RES[15]_2~FF_brt_30_brt_82_brt_151_q ), .I1(\RES[17]_2~FF_brt_8_brt_36_q ), 
            .O(n5129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6821.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6822 (.I0(\RES[15]_2~FF_brt_30_brt_80_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(\RES[15]_2~FF_brt_30_brt_81_q ), .I3(n5129), .O(n5130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__6822.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__6823 (.I0(\RES[15]_2~FF_brt_29_q ), .I1(n5130), .I2(\RES[4]_2~FF_brt_125_q ), 
            .O(n1600_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6823.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6824 (.I0(n3534), .I1(n3527), .I2(\ARG1[31] ), .I3(\SHIFT_STEPS[4] ), 
            .O(n5131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6824.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6825 (.I0(\ARG1[14] ), .I1(\ARG1[16] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6825.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6826 (.I0(n5124), .I1(n5132), .I2(\SHIFT_STEPS[0] ), 
            .O(n5133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6826.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6827 (.I0(n5081), .I1(n5133), .I2(\SHIFT_STEPS[2] ), 
            .O(n5134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6827.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6828 (.I0(n5029), .I1(n5134), .I2(\SHIFT_STEPS[3] ), 
            .I3(n4957), .O(n5135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6828.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6829 (.I0(n5075), .I1(n3542), .I2(n3541), .O(n5136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6829.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6830 (.I0(\RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152_q ), 
            .I1(\RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153_q ), .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), 
            .I3(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .O(n5137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6830.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6831 (.I0(\RES[16]_2~FF_brt_5_brt_33_brt_83_q ), .I1(n5137), 
            .I2(\RES[17]_2~FF_brt_8_brt_36_q ), .O(n5138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6831.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6832 (.I0(\RES[16]_2~FF_brt_5_brt_31_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(\RES[16]_2~FF_brt_5_brt_32_q ), .I3(n5138), .O(n5139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6832.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6833 (.I0(\OPERATION[0] ), .I1(\ARG2[16] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[16] ), .O(n5140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6833.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6834 (.I0(n5131), .I1(n3536), .I2(n5140), .I3(\OPERATION[2] ), 
            .O(n5141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6834.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6835 (.I0(n5139), .I1(\RES[16]_2~FF_brt_6_q ), .I2(\RES[4]_2~FF_brt_125_q ), 
            .O(n1599_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6835.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6836 (.I0(n4969), .I1(n5101), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6836.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6837 (.I0(\ARG1[15] ), .I1(\ARG1[17] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6837.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6838 (.I0(n5132), .I1(n5143), .I2(\SHIFT_STEPS[0] ), 
            .O(n5144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6838.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6839 (.I0(n5043), .I1(n5144), .I2(\SHIFT_STEPS[2] ), 
            .I3(n5142), .O(n5145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6839.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6840 (.I0(\RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154_q ), 
            .I1(\RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155_q ), .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), 
            .I3(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .O(n5146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6840.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6841 (.I0(\RES[17]_2~FF_brt_8_brt_37_brt_85_q ), .I1(\RES[27]_2~FF_brt_53_q ), 
            .I2(\RES[17]_2~FF_brt_8_brt_37_brt_86_q ), .I3(n5146), .O(n5147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__6841.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__6842 (.I0(\RES[17]_2~FF_brt_8_brt_34_q ), .I1(\RES[17]_2~FF_brt_8_brt_35_q ), 
            .I2(\RES[17]_2~FF_brt_8_brt_36_q ), .I3(n5147), .O(n5148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6842.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6843 (.I0(n4886), .I1(n4884), .I2(\SHIFT_STEPS[2] ), 
            .O(n5149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6843.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6844 (.I0(n5149), .I1(n5071), .I2(n5014), .O(n5150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6844.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6845 (.I0(n4881), .I1(n4967), .O(n5151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6845.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6846 (.I0(n5151), .I1(n5150), .I2(n3547), .O(n5152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6846.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6847 (.I0(\OPERATION[0] ), .I1(\ARG2[17] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[17] ), .O(n5153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6847.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6848 (.I0(n5153), .I1(\OPERATION[2] ), .O(n5154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6848.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6849 (.I0(n5151), .I1(n5150), .I2(n3536), .I3(n5154), 
            .O(n5155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6849.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6850 (.I0(\RES[17]_2~FF_brt_7_q ), .I1(n5148), .I2(\RES[17]_2~FF_brt_9_q ), 
            .I3(\RES[4]_2~FF_brt_125_q ), .O(n1598_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6850.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6851 (.I0(n3536), .I1(n5018), .O(n5156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6851.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6852 (.I0(n4923), .I1(\ARG1[31] ), .I2(n5156), .I3(\SHIFT_STEPS[4] ), 
            .O(n5157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__6852.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__6853 (.I0(n5157), .I1(n3552), .O(n5158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6853.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6854 (.I0(n4902), .I1(\SHIFT_STEPS[4] ), .I2(n3542), 
            .I3(\OPERATION[2] ), .O(n5159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__6854.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__6855 (.I0(\ARG1[16] ), .I1(\ARG1[18] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6855.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6856 (.I0(n5143), .I1(n5160), .I2(\SHIFT_STEPS[0] ), 
            .O(n5161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6856.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6857 (.I0(n5107), .I1(n5161), .I2(\SHIFT_STEPS[2] ), 
            .O(n5162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6857.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6858 (.I0(n5056), .I1(n5055), .O(n5163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6858.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6859 (.I0(n5163), .I1(n5162), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__6859.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__6860 (.I0(\OPERATION[0] ), .I1(\OPERATION[1] ), .I2(\ARG2[18] ), 
            .I3(\ARG1[18] ), .O(n5165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd33f */ ;
    defparam LUT__6860.LUTMASK = 16'hd33f;
    EFX_LUT4 LUT__6861 (.I0(\OPERATION[0] ), .I1(\OPERATION[1] ), .I2(\OPERATION[2] ), 
            .O(n5166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6861.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6862 (.I0(n3445), .I1(\ARG2[18] ), .I2(n5166), .I3(n5165), 
            .O(n5167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6862.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6863 (.I0(n5164), .I1(n5159), .I2(n5167), .I3(n5018), 
            .O(n5168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6863.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6864 (.I0(\RES[18]_2~FF_brt_90_brt_156_q ), .I1(\RES[18]_2~FF_brt_90_brt_157_q ), 
            .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .I3(\RES[20]_2~FF_brt_93_brt_164_q ), 
            .O(n5169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6864.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6865 (.I0(\RES[18]_2~FF_brt_88_q ), .I1(\RES[18]_2~FF_brt_89_q ), 
            .I2(n5169), .I3(\RES[4]_2~FF_brt_125_q ), .O(n1597_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6865.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6866 (.I0(n4942), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[4] ), 
            .O(n5170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6866.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6867 (.I0(n5002), .I1(n5065), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6867.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6868 (.I0(\ARG1[17] ), .I1(\ARG1[19] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6868.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6869 (.I0(n5160), .I1(n5172), .I2(\SHIFT_STEPS[0] ), 
            .O(n5173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6869.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6870 (.I0(n5125), .I1(n5173), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n5174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6870.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6871 (.I0(n3542), .I1(\SHIFT_STEPS[4] ), .I2(n4946), 
            .I3(\OPERATION[0] ), .O(n5175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__6871.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__6872 (.I0(n5174), .I1(\SHIFT_STEPS[4] ), .I2(n5171), 
            .I3(n5175), .O(n5176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6872.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6873 (.I0(\OPERATION[2] ), .I1(\OPERATION[1] ), .O(n5177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6873.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6874 (.I0(n5170), .I1(\OPERATION[0] ), .I2(n5176), .I3(n5177), 
            .O(n5178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6874.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6875 (.I0(\OPERATION[0] ), .I1(\ARG2[19] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[19] ), .O(n5179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6875.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6876 (.I0(n5170), .I1(n3536), .I2(n5179), .I3(\OPERATION[2] ), 
            .O(n5180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6876.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6877 (.I0(n1353), .I1(n1412), .I2(\OPERATION[0] ), .I3(n3552), 
            .O(n5181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6877.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6878 (.I0(\RES[19]_2~FF_brt_159_q ), .I1(\RES[19]_2~FF_brt_160_q ), 
            .I2(\RES[19]_2~FF_brt_161_q ), .I3(\RES[4]_2~FF_brt_125_q ), 
            .O(n1596_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6878.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6879 (.I0(n4955), .I1(\ARG1[31] ), .I2(n5156), .I3(\SHIFT_STEPS[4] ), 
            .O(n5182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__6879.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__6880 (.I0(\ARG1[20] ), .I1(\ARG2[20] ), .I2(\OPERATION[0] ), 
            .I3(\OPERATION[2] ), .O(n5183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__6880.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__6881 (.I0(\ARG2[20] ), .I1(\ARG1[20] ), .I2(n5183), 
            .I3(\OPERATION[1] ), .O(n5184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ff0 */ ;
    defparam LUT__6881.LUTMASK = 16'h1ff0;
    EFX_LUT4 LUT__6882 (.I0(n5182), .I1(n5184), .O(n5185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6882.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6883 (.I0(\ARG1[18] ), .I1(\ARG1[20] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6883.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6884 (.I0(n5172), .I1(n5186), .I2(\SHIFT_STEPS[0] ), 
            .O(n5187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6884.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6885 (.I0(n5133), .I1(n5187), .I2(\SHIFT_STEPS[2] ), 
            .O(n5188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6885.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6886 (.I0(n5082), .I1(n5188), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6886.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6887 (.I0(n4961), .I1(n5005), .I2(n5189), .I3(n5000), 
            .O(n5190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6887.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6888 (.I0(\RES[20]_2~FF_brt_93_brt_162_q ), .I1(\RES[20]_2~FF_brt_93_brt_163_q ), 
            .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .I3(\RES[20]_2~FF_brt_93_brt_164_q ), 
            .O(n5191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6888.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6889 (.I0(\RES[20]_2~FF_brt_91_q ), .I1(\RES[20]_2~FF_brt_92_q ), 
            .I2(n5191), .I3(\RES[4]_2~FF_brt_125_q ), .O(n1595_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6889.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6890 (.I0(n4978), .I1(\ARG1[31] ), .I2(n5156), .I3(\SHIFT_STEPS[4] ), 
            .O(n5192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__6890.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__6891 (.I0(n5102), .I1(n5071), .I2(n5177), .O(n5193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6891.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6892 (.I0(\ARG1[19] ), .I1(\ARG1[21] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6892.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6893 (.I0(n5186), .I1(n5194), .I2(\SHIFT_STEPS[0] ), 
            .O(n5195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6893.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6894 (.I0(n5144), .I1(n5195), .I2(\SHIFT_STEPS[2] ), 
            .O(n5196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6894.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6895 (.I0(n4970), .I1(n5196), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[4] ), .O(n5197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6895.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6896 (.I0(\OPERATION[0] ), .I1(\ARG2[21] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[21] ), .O(n5198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6896.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6897 (.I0(n3547), .I1(n5198), .I2(\OPERATION[2] ), .O(n5199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6897.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6898 (.I0(n5197), .I1(n5193), .I2(n5199), .O(n5200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6898.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6899 (.I0(\RES[21]_2~FF_brt_96_brt_165_q ), .I1(\RES[21]_2~FF_brt_96_brt_166_q ), 
            .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .I3(\RES[20]_2~FF_brt_93_brt_164_q ), 
            .O(n5201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6899.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6900 (.I0(\RES[21]_2~FF_brt_94_q ), .I1(\RES[21]_2~FF_brt_95_q ), 
            .I2(n5201), .I3(\RES[4]_2~FF_brt_125_q ), .O(n1594_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__6900.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__6901 (.I0(\RES[22]_2~FF_brt_41_brt_97_brt_167_q ), .I1(\RES[22]_2~FF_brt_41_brt_97_brt_168_q ), 
            .I2(\RES[22]_2~FF_brt_41_brt_97_brt_169_q ), .O(n5202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6901.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6902 (.I0(n5202), .I1(\RES[20]_2~FF_brt_93_brt_164_q ), 
            .I2(\RES[22]_2~FF_brt_41_brt_98_q ), .O(n5203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6902.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6903 (.I0(n4990), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[4] ), 
            .O(n5204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6903.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6904 (.I0(\OPERATION[0] ), .I1(\ARG2[22] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[22] ), .O(n5205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6904.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6905 (.I0(n5166), .I1(n5205), .O(n5206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6905.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6906 (.I0(n5086), .I1(n3536), .I2(n5206), .I3(n5204), 
            .O(n5207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa30 */ ;
    defparam LUT__6906.LUTMASK = 16'hfa30;
    EFX_LUT4 LUT__6907 (.I0(\ARG1[20] ), .I1(\ARG1[22] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6907.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6908 (.I0(n5194), .I1(n5208), .I2(\SHIFT_STEPS[0] ), 
            .O(n5209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6908.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6909 (.I0(n5161), .I1(n5209), .I2(\SHIFT_STEPS[2] ), 
            .O(n5210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6909.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6910 (.I0(n5109), .I1(n5210), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6910.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6911 (.I0(n4994), .I1(n5005), .I2(n5211), .I3(n5000), 
            .O(n5212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__6911.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__6912 (.I0(\RES[22]_2~FF_brt_38_q ), .I1(\RES[22]_2~FF_brt_39_q ), 
            .I2(\RES[20]_2~FF_brt_93_brt_164_q ), .I3(n5203), .O(n1593_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__6912.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__6913 (.I0(n5008), .I1(\ARG1[31] ), .I2(n5156), .I3(n4967), 
            .O(n5213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__6913.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__6914 (.I0(\ARG1[21] ), .I1(\ARG1[23] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6914.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6915 (.I0(n5208), .I1(n5214), .I2(\SHIFT_STEPS[0] ), 
            .O(n5215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6915.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6916 (.I0(n5173), .I1(n5215), .I2(\SHIFT_STEPS[2] ), 
            .O(n5216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6916.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6917 (.I0(n5126), .I1(n5216), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6917.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6918 (.I0(n5003), .I1(n5005), .I2(n5217), .I3(n5000), 
            .O(n5218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6918.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6919 (.I0(\OPERATION[0] ), .I1(\ARG2[23] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[23] ), .O(n5219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6919.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6920 (.I0(\OPERATION[1] ), .I1(n5219), .I2(\OPERATION[2] ), 
            .O(n5220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6920.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6921 (.I0(\RES[23]_2~FF_brt_45_brt_99_brt_170_q ), .I1(\RES[23]_2~FF_brt_45_brt_99_brt_171_q ), 
            .I2(\RES[22]_2~FF_brt_41_brt_97_brt_169_q ), .O(n5221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6921.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6922 (.I0(n5221), .I1(\RES[23]_2~FF_brt_45_brt_100_q ), 
            .I2(\RES[4]_2~FF_brt_125_q ), .O(n5222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6922.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6923 (.I0(\RES[23]_2~FF_brt_42_q ), .I1(\RES[23]_2~FF_brt_43_q ), 
            .I2(\RES[23]_2~FF_brt_44_q ), .I3(n5222), .O(n1592_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6923.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6924 (.I0(n3526), .I1(n3523), .I2(\SHIFT_STEPS[2] ), 
            .O(n5223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6924.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6925 (.I0(n5223), .I1(\ARG1[31] ), .I2(n4967), .I3(n3536), 
            .O(n5224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6925.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6926 (.I0(\OPERATION[0] ), .I1(\ARG2[24] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[24] ), .O(n5225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6926.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6927 (.I0(\ARG1[22] ), .I1(\ARG1[24] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6927.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6928 (.I0(n5214), .I1(n5226), .I2(\SHIFT_STEPS[0] ), 
            .O(n5227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6928.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6929 (.I0(n5187), .I1(n5227), .I2(\SHIFT_STEPS[2] ), 
            .O(n5228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6929.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6930 (.I0(n5134), .I1(n5228), .I2(\SHIFT_STEPS[3] ), 
            .I3(n4957), .O(n5229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__6930.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__6931 (.I0(n5029), .I1(\SHIFT_STEPS[3] ), .I2(n5031), 
            .I3(n5075), .O(n5230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__6931.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__6932 (.I0(n5223), .I1(\ARG1[31] ), .I2(n4967), .I3(n3547), 
            .O(n5231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__6932.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__6933 (.I0(\OPERATION[1] ), .I1(\OPERATION[0] ), .O(n5232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6933.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6934 (.I0(n3536), .I1(n1402), .I2(n3545), .O(n5233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__6934.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__6935 (.I0(\RES[24]_2~FF_brt_49_brt_105_brt_172_q ), .I1(\RES[24]_2~FF_brt_49_brt_105_brt_173_q ), 
            .I2(\RES[24]_2~FF_brt_49_brt_105_brt_174_q ), .O(n5234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__6935.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__6936 (.I0(\RES[24]_2~FF_brt_49_brt_102_q ), .I1(\RES[24]_2~FF_brt_49_brt_103_q ), 
            .I2(\RES[24]_2~FF_brt_49_brt_104_q ), .I3(n5234), .O(n5235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6936.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6937 (.I0(\RES[24]_2~FF_brt_46_q ), .I1(\RES[24]_2~FF_brt_47_q ), 
            .I2(\RES[24]_2~FF_brt_48_q ), .I3(n5235), .O(n1591_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__6937.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__6938 (.I0(\ARG1[23] ), .I1(\ARG1[25] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6938.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6939 (.I0(n5226), .I1(n5236), .I2(\SHIFT_STEPS[0] ), 
            .O(n5237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6939.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6940 (.I0(n5195), .I1(n5237), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n5238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6940.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6941 (.I0(n5101), .I1(n5144), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6941.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6942 (.I0(n5239), .I1(n5238), .I2(n4957), .O(n5240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6942.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6943 (.I0(n5044), .I1(\SHIFT_STEPS[3] ), .I2(n5045), 
            .I3(n5075), .O(n5241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__6943.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__6944 (.I0(n5149), .I1(\ARG1[31] ), .I2(n4967), .I3(n3547), 
            .O(n5242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6944.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6945 (.I0(n3536), .I1(n1400), .I2(n3545), .O(n5243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__6945.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__6946 (.I0(\RES[24]_2~FF_brt_49_brt_105_brt_172_q ), .I1(\RES[25]_2~FF_brt_108_brt_175_q ), 
            .I2(\RES[25]_2~FF_brt_108_brt_176_q ), .I3(\RES[25]_2~FF_brt_108_brt_177_q ), 
            .O(n5244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6946.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6947 (.I0(\OPERATION[0] ), .I1(\ARG2[25] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[25] ), .O(n5245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6947.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6948 (.I0(n5149), .I1(\ARG1[31] ), .I2(n4967), .I3(n3536), 
            .O(n5246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6948.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6949 (.I0(n5246), .I1(n5245), .I2(n3537), .O(n5247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6949.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6950 (.I0(\RES[25]_2~FF_brt_106_q ), .I1(\RES[25]_2~FF_brt_107_q ), 
            .I2(n5244), .I3(\RES[25]_2~FF_brt_109_q ), .O(n1590_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__6950.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__6951 (.I0(n5058), .I1(n5075), .O(n5248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6951.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6952 (.I0(n4922), .I1(\ARG1[31] ), .I2(n4967), .O(n5249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6952.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6953 (.I0(\ARG1[24] ), .I1(\ARG1[26] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6953.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6954 (.I0(n5236), .I1(n5250), .I2(\SHIFT_STEPS[0] ), 
            .O(n5251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6954.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6955 (.I0(n5209), .I1(n5251), .I2(\SHIFT_STEPS[2] ), 
            .O(n5252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6955.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6956 (.I0(n5162), .I1(n5252), .I2(\SHIFT_STEPS[3] ), 
            .I3(n4957), .O(n5253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6956.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6957 (.I0(\RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178_q ), 
            .I1(\RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179_q ), .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), 
            .I3(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .O(n5254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6957.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6958 (.I0(n5254), .I1(\RES[17]_2~FF_brt_8_brt_36_q ), 
            .O(n5255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6958.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6959 (.I0(\RES[26]_2~FF_brt_10_brt_50_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(\RES[26]_2~FF_brt_10_brt_51_q ), .I3(n5255), .O(n5256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__6959.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__6960 (.I0(\OPERATION[0] ), .I1(\ARG2[26] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[26] ), .O(n5257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6960.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6961 (.I0(n5249), .I1(n3536), .I2(n5257), .I3(\OPERATION[2] ), 
            .O(n5258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6961.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6962 (.I0(n5256), .I1(\RES[26]_2~FF_brt_11_q ), .I2(\RES[26]_2~FF_brt_12_q ), 
            .I3(\RES[4]_2~FF_brt_125_q ), .O(n1589_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__6962.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__6963 (.I0(n5125), .I1(n5173), .I2(\SHIFT_STEPS[2] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6963.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6964 (.I0(\ARG1[25] ), .I1(\ARG1[27] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6964.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6965 (.I0(n5250), .I1(n5260), .I2(\SHIFT_STEPS[0] ), 
            .O(n5261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6965.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6966 (.I0(n5215), .I1(n5261), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[2] ), .O(n5262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6966.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6967 (.I0(n5007), .I1(\ARG1[31] ), .I2(n4903), .O(n5263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__6967.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__6968 (.I0(n1345), .I1(n1396), .I2(\OPERATION[1] ), .I3(\OPERATION[0] ), 
            .O(n5264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6968.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6969 (.I0(\RES[27]_2~FF_brt_55_brt_113_brt_180_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(\RES[27]_2~FF_brt_55_brt_113_brt_181_q ), .I3(\RES[28]_2~FF_brt_14_q ), 
            .O(n5265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__6969.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__6970 (.I0(\RES[27]_2~FF_brt_55_brt_111_q ), .I1(\RES[27]_2~FF_brt_55_brt_112_q ), 
            .I2(\RES[17]_2~FF_brt_8_brt_34_q ), .I3(n5265), .O(n5266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6970.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6971 (.I0(\OPERATION[0] ), .I1(\ARG1[27] ), .I2(\OPERATION[1] ), 
            .I3(\ARG2[27] ), .O(n5267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6971.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6972 (.I0(n3536), .I1(n5263), .I2(n5267), .I3(n3537), 
            .O(n5268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6972.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6973 (.I0(\RES[27]_2~FF_brt_53_q ), .I1(\RES[27]_2~FF_brt_54_q ), 
            .I2(n5266), .I3(\RES[27]_2~FF_brt_56_q ), .O(n1588_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__6973.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__6974 (.I0(n3523), .I1(\ARG1[31] ), .I2(n4903), .O(n5269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__6974.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__6975 (.I0(\OPERATION[0] ), .I1(\ARG1[28] ), .I2(\OPERATION[1] ), 
            .I3(\ARG2[28] ), .O(n5270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6975.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6976 (.I0(n3536), .I1(n5269), .I2(n5270), .I3(\OPERATION[3] ), 
            .O(n5271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__6976.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__6977 (.I0(\ARG1[26] ), .I1(\ARG1[28] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6977.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6978 (.I0(n5272), .I1(n5260), .I2(\SHIFT_STEPS[0] ), 
            .O(n5273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6978.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6979 (.I0(n5227), .I1(n5273), .I2(\SHIFT_STEPS[2] ), 
            .O(n5274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6979.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6980 (.I0(n5188), .I1(n5274), .I2(\SHIFT_STEPS[4] ), 
            .I3(\SHIFT_STEPS[3] ), .O(n5275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__6980.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__6981 (.I0(n4961), .I1(n5082), .I2(\SHIFT_STEPS[3] ), 
            .I3(\SHIFT_STEPS[4] ), .O(n5276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6981.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6982 (.I0(\RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182_q ), 
            .I1(\RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_q ), .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), 
            .I3(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .O(n5277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6982.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6983 (.I0(\RES[28]_2~FF_brt_15_brt_60_brt_114_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(n5277), .I3(\RES[17]_2~FF_brt_8_brt_36_q ), .O(n5278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6983.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6984 (.I0(\RES[28]_2~FF_brt_15_brt_57_q ), .I1(\RES[28]_2~FF_brt_15_brt_58_q ), 
            .I2(\RES[28]_2~FF_brt_15_brt_59_q ), .I3(n5278), .O(n5279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6984.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6985 (.I0(\RES[28]_2~FF_brt_13_q ), .I1(\RES[28]_2~FF_brt_14_q ), 
            .I2(n5279), .O(n1587_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6985.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6986 (.I0(\ARG1[27] ), .I1(\ARG1[29] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6986.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6987 (.I0(n5272), .I1(n5280), .I2(\SHIFT_STEPS[0] ), 
            .O(n5281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6987.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6988 (.I0(n5237), .I1(n5281), .I2(\SHIFT_STEPS[2] ), 
            .O(n5282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__6988.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__6989 (.I0(n5196), .I1(n5282), .I2(\SHIFT_STEPS[3] ), 
            .I3(n4957), .O(n5283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6989.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6990 (.I0(n4977), .I1(\ARG1[31] ), .I2(n4967), .O(n5284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6990.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6991 (.I0(\RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184_q ), 
            .I1(\RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185_q ), .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), 
            .I3(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_138_q ), .O(n5285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6991.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6992 (.I0(\RES[29]_2~FF_brt_16_brt_63_brt_116_q ), .I1(\RES[9]_2~FF_brt_1_brt_24_q ), 
            .I2(n5285), .I3(\RES[17]_2~FF_brt_8_brt_36_q ), .O(n5286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6992.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6993 (.I0(\RES[29]_2~FF_brt_16_brt_61_q ), .I1(\RES[27]_2~FF_brt_53_q ), 
            .I2(\RES[29]_2~FF_brt_16_brt_62_q ), .I3(n5286), .O(n5287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6993.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6994 (.I0(\OPERATION[0] ), .I1(\ARG1[29] ), .I2(\OPERATION[1] ), 
            .I3(\ARG2[29] ), .O(n5288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__6994.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__6995 (.I0(n5284), .I1(n3536), .I2(n5288), .I3(\OPERATION[2] ), 
            .O(n5289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6995.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6996 (.I0(n5287), .I1(\RES[29]_2~FF_brt_17_q ), .I2(\RES[4]_2~FF_brt_125_q ), 
            .O(n1586_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6996.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6997 (.I0(\ARG1[28] ), .I1(\ARG1[30] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__6997.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__6998 (.I0(n5280), .I1(n5290), .I2(\SHIFT_STEPS[0] ), 
            .O(n5291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6998.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6999 (.I0(n5251), .I1(n5291), .I2(\SHIFT_STEPS[2] ), 
            .O(n5292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__6999.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__7000 (.I0(n5210), .I1(n5292), .I2(\SHIFT_STEPS[3] ), 
            .O(n5293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7000.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7001 (.I0(n5110), .I1(n5293), .I2(\SHIFT_STEPS[4] ), 
            .I3(n3445), .O(n5294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__7001.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__7002 (.I0(n1390), .I1(n1342), .I2(\OPERATION[1] ), .I3(n5166), 
            .O(n5295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7002.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7003 (.I0(n4921), .I1(\ARG1[31] ), .I2(n4903), .O(n5296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__7003.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__7004 (.I0(n5296), .I1(n3547), .I2(n3545), .O(n5297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__7004.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__7005 (.I0(\OPERATION[0] ), .I1(\ARG2[30] ), .I2(\OPERATION[1] ), 
            .I3(\ARG1[30] ), .O(n5298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h873f */ ;
    defparam LUT__7005.LUTMASK = 16'h873f;
    EFX_LUT4 LUT__7006 (.I0(n3536), .I1(n5296), .I2(n5298), .I3(n3537), 
            .O(n5299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__7006.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__7007 (.I0(\RES[30]_2~FF_brt_186_q ), .I1(\RES[30]_2~FF_brt_187_q ), 
            .I2(\RES[30]_2~FF_brt_188_q ), .I3(\RES[30]_2~FF_brt_189_q ), 
            .O(n1585_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__7007.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__7008 (.I0(n5003), .I1(n5126), .I2(\SHIFT_STEPS[3] ), 
            .I3(n5075), .O(n5300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7008.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7009 (.I0(\ARG1[29] ), .I1(\ARG1[31] ), .I2(\SHIFT_STEPS[1] ), 
            .O(n5301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7009.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7010 (.I0(n5290), .I1(n5301), .I2(\SHIFT_STEPS[0] ), 
            .O(n5302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7010.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7011 (.I0(n5261), .I1(n5302), .I2(\SHIFT_STEPS[2] ), 
            .O(n5303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7011.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7012 (.I0(n5216), .I1(n5303), .I2(\SHIFT_STEPS[3] ), 
            .I3(n4957), .O(n5304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__7012.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__7013 (.I0(\RES[31]_2~FF_brt_66_brt_119_brt_190_q ), .I1(\RES[31]_2~FF_brt_66_brt_119_brt_191_q ), 
            .I2(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q ), .I3(\RES[22]_2~FF_brt_41_brt_97_brt_169_q ), 
            .O(n5305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__7013.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__7014 (.I0(\RES[9]_2~FF_brt_1_brt_24_q ), .I1(\RES[31]_2~FF_brt_66_brt_118_q ), 
            .I2(\RES[17]_2~FF_brt_8_brt_36_q ), .I3(n5305), .O(n5306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__7014.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__7015 (.I0(\OPERATION[0] ), .I1(\ARG1[31] ), .I2(\OPERATION[1] ), 
            .I3(\ARG2[31] ), .O(n5307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h833b */ ;
    defparam LUT__7015.LUTMASK = 16'h833b;
    EFX_LUT4 LUT__7016 (.I0(n5307), .I1(\OPERATION[2] ), .I2(\OPERATION[3] ), 
            .O(n5308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__7016.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__7017 (.I0(\RES[31]_2~FF_brt_64_q ), .I1(\RES[31]_2~FF_brt_65_q ), 
            .I2(n5306), .I3(\RES[31]_2~FF_brt_67_q ), .O(n1584_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__7017.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__7018 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[8] ), .O(n1575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7018.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7019 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[9] ), .O(n1574_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7019.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7020 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[10] ), .O(n1573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7020.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7021 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[11] ), .O(n1572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7021.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7022 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[12] ), .O(n1571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7022.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7023 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[13] ), .O(n1570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7023.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7024 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[14] ), .O(n1569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7024.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7025 (.I0(\DATA_FORMAT_2[2] ), .I1(\ARG2[15] ), .O(n1568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7025.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7026 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[16] ), .O(n1567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7026.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7027 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[17] ), .O(n1566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7027.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7028 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[18] ), .O(n1565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7028.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7029 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[19] ), .O(n1564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7029.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7030 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[20] ), .O(n1563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7030.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7031 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[21] ), .O(n1562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7031.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7032 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[22] ), .O(n1561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7032.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7033 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[23] ), .O(n1560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7033.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7034 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[24] ), .O(n1559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7034.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7035 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[25] ), .O(n1558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7035.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7036 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[26] ), .O(n1557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7036.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7037 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[27] ), .O(n1556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7037.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7038 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[28] ), .O(n1555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7038.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7039 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[29] ), .O(n1554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7039.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7040 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[30] ), .O(n1553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7040.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7041 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[2] ), 
            .I2(\ARG2[31] ), .O(n1552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7041.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7042 (.I0(\LOAD_DATA[8] ), .I1(\XI[0][8] ), .I2(n4733), 
            .O(n5309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7042.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7043 (.I0(\DATA_FORMAT_2[2] ), .I1(LOAD_OP), .O(n5310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7043.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7044 (.I0(n5310), .I1(\DATA_FORMAT_2[0] ), .O(n5311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7044.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7045 (.I0(\DATA_FORMAT_2[0] ), .I1(\DATA_FORMAT_2[1] ), 
            .I2(\DATA_FORMAT_2[2] ), .I3(LOAD_OP), .O(n5312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__7045.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__7046 (.I0(\LOAD_DATA[7] ), .I1(\DATA_FORMAT_2[2] ), .I2(n5312), 
            .O(n5313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7046.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7047 (.I0(n5309), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7047.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7048 (.I0(n5309), .I1(n5311), .I2(n5313), .I3(n5314), 
            .O(n17577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7048.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7049 (.I0(\DATA_FORMAT_2[2] ), .I1(\DATA_FORMAT_2[1] ), 
            .I2(\DATA_FORMAT_2[0] ), .I3(LOAD_OP), .O(n5315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__7049.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__7050 (.I0(n4733), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net41512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7050.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7051 (.I0(\LOAD_DATA[9] ), .I1(\XI[0][9] ), .I2(n4733), 
            .O(n5316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7051.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7052 (.I0(n5316), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7052.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7053 (.I0(n5316), .I1(n5311), .I2(n5313), .I3(n5317), 
            .O(n17576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7053.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7054 (.I0(\LOAD_DATA[10] ), .I1(\XI[0][10] ), .I2(n4733), 
            .O(n5318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7054.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7055 (.I0(n5318), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7055.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7056 (.I0(n5318), .I1(n5311), .I2(n5313), .I3(n5319), 
            .O(n17575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7056.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7057 (.I0(\LOAD_DATA[11] ), .I1(\XI[0][11] ), .I2(n4733), 
            .O(n5320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7057.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7058 (.I0(n5320), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7058.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7059 (.I0(n5320), .I1(n5311), .I2(n5313), .I3(n5321), 
            .O(n17574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7059.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7060 (.I0(\LOAD_DATA[12] ), .I1(\XI[0][12] ), .I2(n4733), 
            .O(n5322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7060.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7061 (.I0(n5322), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7061.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7062 (.I0(n5322), .I1(n5311), .I2(n5313), .I3(n5323), 
            .O(n17573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7062.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7063 (.I0(\LOAD_DATA[13] ), .I1(\XI[0][13] ), .I2(n4733), 
            .O(n5324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7063.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7064 (.I0(n5324), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7064.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7065 (.I0(n5324), .I1(n5311), .I2(n5313), .I3(n5325), 
            .O(n17572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7065.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7066 (.I0(\LOAD_DATA[14] ), .I1(\XI[0][14] ), .I2(n4733), 
            .O(n5326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7066.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7067 (.I0(n5326), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7067.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7068 (.I0(n5326), .I1(n5311), .I2(n5313), .I3(n5327), 
            .O(n17571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7068.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7069 (.I0(\LOAD_DATA[15] ), .I1(\XI[0][15] ), .I2(n4733), 
            .O(n5328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7069.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7070 (.I0(n5328), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7070.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7071 (.I0(n5328), .I1(n5311), .I2(n5313), .I3(n5329), 
            .O(n17570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7071.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7072 (.I0(\DATA_FORMAT_2[1] ), .I1(\LOAD_DATA[15] ), .I2(\DATA_FORMAT_2[0] ), 
            .I3(\DATA_FORMAT_2[2] ), .O(n5330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__7072.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__7073 (.I0(n4733), .I1(n5330), .O(n5331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7073.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7074 (.I0(\DATA_FORMAT_2[0] ), .I1(\LOAD_DATA[7] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[2] ), .O(n5332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7074.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7075 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[16] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7075.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7076 (.I0(n5333), .I1(n5332), .I2(LOAD_OP), .O(n5334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__7076.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__7077 (.I0(LOAD_OP), .I1(n1599_2), .O(n5335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7077.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7078 (.I0(\XI[0][16] ), .I1(n5331), .I2(n5334), .I3(n5335), 
            .O(n17569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7078.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7079 (.I0(\DATA_FORMAT_2[1] ), .I1(\DATA_FORMAT_2[0] ), 
            .I2(\DATA_FORMAT_2[2] ), .I3(LOAD_OP), .O(n5336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__7079.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__7080 (.I0(n4733), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net49709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7080.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7081 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[17] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7081.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7082 (.I0(n5332), .I1(n5337), .I2(LOAD_OP), .O(n5338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7082.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7083 (.I0(LOAD_OP), .I1(n1598_2), .O(n5339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7083.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7084 (.I0(\XI[0][17] ), .I1(n5331), .I2(n5338), .I3(n5339), 
            .O(n17568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7084.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7085 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[18] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7085.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7086 (.I0(n5332), .I1(n5340), .I2(LOAD_OP), .O(n5341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7086.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7087 (.I0(LOAD_OP), .I1(n1597_2), .O(n5342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7087.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7088 (.I0(\XI[0][18] ), .I1(n5331), .I2(n5341), .I3(n5342), 
            .O(n17567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7088.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7089 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[19] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7089.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7090 (.I0(n5332), .I1(n5343), .I2(LOAD_OP), .O(n5344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7090.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7091 (.I0(LOAD_OP), .I1(n1596_2), .O(n5345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7091.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7092 (.I0(\XI[0][19] ), .I1(n5331), .I2(n5344), .I3(n5345), 
            .O(n17566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7092.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7093 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[20] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7093.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7094 (.I0(n5332), .I1(n5346), .I2(LOAD_OP), .O(n5347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7094.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7095 (.I0(LOAD_OP), .I1(n1595_2), .O(n5348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7095.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7096 (.I0(\XI[0][20] ), .I1(n5331), .I2(n5347), .I3(n5348), 
            .O(n17565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7096.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7097 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[21] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7097.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7098 (.I0(n5332), .I1(n5349), .I2(LOAD_OP), .O(n5350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7098.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7099 (.I0(LOAD_OP), .I1(n1594_2), .O(n5351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7099.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7100 (.I0(\XI[0][21] ), .I1(n5331), .I2(n5350), .I3(n5351), 
            .O(n17564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7100.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7101 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[22] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7101.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7102 (.I0(n5332), .I1(n5352), .I2(LOAD_OP), .O(n5353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7102.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7103 (.I0(LOAD_OP), .I1(n1593_2), .O(n5354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7103.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7104 (.I0(\XI[0][22] ), .I1(n5331), .I2(n5353), .I3(n5354), 
            .O(n17563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7104.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7105 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[23] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7105.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7106 (.I0(n5332), .I1(n5355), .I2(LOAD_OP), .O(n5356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7106.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7107 (.I0(LOAD_OP), .I1(n1592_2), .O(n5357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7107.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7108 (.I0(\XI[0][23] ), .I1(n5331), .I2(n5356), .I3(n5357), 
            .O(n17562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7108.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7109 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[24] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7109.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7110 (.I0(n5332), .I1(n5358), .I2(LOAD_OP), .O(n5359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7110.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7111 (.I0(LOAD_OP), .I1(n1591_2), .O(n5360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7111.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7112 (.I0(\XI[0][24] ), .I1(n5331), .I2(n5359), .I3(n5360), 
            .O(n17561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7112.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7113 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[25] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7113.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7114 (.I0(n5332), .I1(n5361), .I2(LOAD_OP), .O(n5362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7114.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7115 (.I0(LOAD_OP), .I1(n1590_2), .O(n5363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7115.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7116 (.I0(\XI[0][25] ), .I1(n5331), .I2(n5362), .I3(n5363), 
            .O(n17560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7116.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7117 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[26] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7117.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7118 (.I0(n5332), .I1(n5364), .I2(LOAD_OP), .O(n5365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7118.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7119 (.I0(LOAD_OP), .I1(n1589_2), .O(n5366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7119.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7120 (.I0(\XI[0][26] ), .I1(n5331), .I2(n5365), .I3(n5366), 
            .O(n17559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7120.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7121 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[27] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7121.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7122 (.I0(n5332), .I1(n5367), .I2(LOAD_OP), .O(n5368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7122.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7123 (.I0(LOAD_OP), .I1(n1588_2), .O(n5369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7123.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7124 (.I0(\XI[0][27] ), .I1(n5331), .I2(n5368), .I3(n5369), 
            .O(n17558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7124.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7125 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[28] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7125.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7126 (.I0(n5332), .I1(n5370), .I2(LOAD_OP), .O(n5371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7126.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7127 (.I0(LOAD_OP), .I1(n1587_2), .O(n5372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7127.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7128 (.I0(\XI[0][28] ), .I1(n5331), .I2(n5371), .I3(n5372), 
            .O(n17557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7128.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7129 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[29] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7129.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7130 (.I0(n5332), .I1(n5373), .I2(LOAD_OP), .O(n5374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7130.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7131 (.I0(LOAD_OP), .I1(n1586_2), .O(n5375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7131.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7132 (.I0(\XI[0][29] ), .I1(n5331), .I2(n5374), .I3(n5375), 
            .O(n17556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7132.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7133 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[30] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7133.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7134 (.I0(n5332), .I1(n5376), .I2(LOAD_OP), .O(n5377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7134.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7135 (.I0(LOAD_OP), .I1(n1585_2), .O(n5378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7135.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7136 (.I0(\XI[0][30] ), .I1(n5331), .I2(n5377), .I3(n5378), 
            .O(n17555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7136.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7137 (.I0(\LOAD_DATA[15] ), .I1(\LOAD_DATA[31] ), .I2(\DATA_FORMAT_2[1] ), 
            .I3(\DATA_FORMAT_2[0] ), .O(n5379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7137.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7138 (.I0(n5332), .I1(n5379), .I2(LOAD_OP), .O(n5380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7138.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7139 (.I0(LOAD_OP), .I1(n1584_2), .O(n5381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7139.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7140 (.I0(\XI[0][31] ), .I1(n5331), .I2(n5380), .I3(n5381), 
            .O(n17554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7140.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7141 (.I0(\LOAD_DATA[8] ), .I1(\XI[1][8] ), .I2(n4735), 
            .O(n5382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7141.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7142 (.I0(n5382), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7142.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7143 (.I0(n5382), .I1(n5311), .I2(n5313), .I3(n5383), 
            .O(n17610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7143.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7144 (.I0(n4735), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net41704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7144.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7145 (.I0(\LOAD_DATA[9] ), .I1(\XI[1][9] ), .I2(n4735), 
            .O(n5384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7145.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7146 (.I0(n5384), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7146.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7147 (.I0(n5384), .I1(n5311), .I2(n5313), .I3(n5385), 
            .O(n17609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7147.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7148 (.I0(\LOAD_DATA[10] ), .I1(\XI[1][10] ), .I2(n4735), 
            .O(n5386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7148.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7149 (.I0(n5386), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7149.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7150 (.I0(n5386), .I1(n5311), .I2(n5313), .I3(n5387), 
            .O(n17608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7150.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7151 (.I0(\LOAD_DATA[11] ), .I1(\XI[1][11] ), .I2(n4735), 
            .O(n5388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7151.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7152 (.I0(n5388), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7152.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7153 (.I0(n5388), .I1(n5311), .I2(n5313), .I3(n5389), 
            .O(n17607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7153.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7154 (.I0(\LOAD_DATA[12] ), .I1(\XI[1][12] ), .I2(n4735), 
            .O(n5390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7154.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7155 (.I0(n5390), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7155.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7156 (.I0(n5390), .I1(n5311), .I2(n5313), .I3(n5391), 
            .O(n17606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7156.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7157 (.I0(\LOAD_DATA[13] ), .I1(\XI[1][13] ), .I2(n4735), 
            .O(n5392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7157.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7158 (.I0(n5392), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7158.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7159 (.I0(n5392), .I1(n5311), .I2(n5313), .I3(n5393), 
            .O(n17605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7159.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7160 (.I0(\LOAD_DATA[14] ), .I1(\XI[1][14] ), .I2(n4735), 
            .O(n5394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7160.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7161 (.I0(n5394), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7161.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7162 (.I0(n5394), .I1(n5311), .I2(n5313), .I3(n5395), 
            .O(n17604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7162.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7163 (.I0(\LOAD_DATA[15] ), .I1(\XI[1][15] ), .I2(n4735), 
            .O(n5396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7163.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7164 (.I0(n5396), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7164.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7165 (.I0(n5396), .I1(n5311), .I2(n5313), .I3(n5397), 
            .O(n17603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7165.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7166 (.I0(n4735), .I1(n5330), .O(n5398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7166.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7167 (.I0(\XI[1][16] ), .I1(n5398), .I2(n5334), .I3(n5335), 
            .O(n17602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7167.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7168 (.I0(n4735), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net49773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7168.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7169 (.I0(\XI[1][17] ), .I1(n5398), .I2(n5338), .I3(n5339), 
            .O(n17601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7169.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7170 (.I0(\XI[1][18] ), .I1(n5398), .I2(n5341), .I3(n5342), 
            .O(n17600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7170.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7171 (.I0(\XI[1][19] ), .I1(n5398), .I2(n5344), .I3(n5345), 
            .O(n17599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7171.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7172 (.I0(\XI[1][20] ), .I1(n5398), .I2(n5347), .I3(n5348), 
            .O(n17598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7172.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7173 (.I0(\XI[1][21] ), .I1(n5398), .I2(n5350), .I3(n5351), 
            .O(n17597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7173.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7174 (.I0(\XI[1][22] ), .I1(n5398), .I2(n5353), .I3(n5354), 
            .O(n17596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7174.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7175 (.I0(\XI[1][23] ), .I1(n5398), .I2(n5356), .I3(n5357), 
            .O(n17595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7175.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7176 (.I0(\XI[1][24] ), .I1(n5398), .I2(n5359), .I3(n5360), 
            .O(n17594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7176.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7177 (.I0(\XI[1][25] ), .I1(n5398), .I2(n5362), .I3(n5363), 
            .O(n17593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7177.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7178 (.I0(\XI[1][26] ), .I1(n5398), .I2(n5365), .I3(n5366), 
            .O(n17592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7178.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7179 (.I0(\XI[1][27] ), .I1(n5398), .I2(n5368), .I3(n5369), 
            .O(n17591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7179.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7180 (.I0(\XI[1][28] ), .I1(n5398), .I2(n5371), .I3(n5372), 
            .O(n17590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7180.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7181 (.I0(\XI[1][29] ), .I1(n5398), .I2(n5374), .I3(n5375), 
            .O(n17589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7181.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7182 (.I0(\XI[1][30] ), .I1(n5398), .I2(n5377), .I3(n5378), 
            .O(n17588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7182.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7183 (.I0(\XI[1][31] ), .I1(n5398), .I2(n5380), .I3(n5381), 
            .O(n17587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7183.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7184 (.I0(\LOAD_DATA[8] ), .I1(\XI[2][8] ), .I2(n4737), 
            .O(n5399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7184.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7185 (.I0(n5399), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7185.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7186 (.I0(n5399), .I1(n5311), .I2(n5313), .I3(n5400), 
            .O(n17643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7186.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7187 (.I0(n4737), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net41896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7187.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7188 (.I0(\LOAD_DATA[9] ), .I1(\XI[2][9] ), .I2(n4737), 
            .O(n5401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7188.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7189 (.I0(n5401), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7189.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7190 (.I0(n5401), .I1(n5311), .I2(n5313), .I3(n5402), 
            .O(n17642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7190.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7191 (.I0(\LOAD_DATA[10] ), .I1(\XI[2][10] ), .I2(n4737), 
            .O(n5403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7191.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7192 (.I0(n5403), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7192.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7193 (.I0(n5403), .I1(n5311), .I2(n5313), .I3(n5404), 
            .O(n17641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7193.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7194 (.I0(\LOAD_DATA[11] ), .I1(\XI[2][11] ), .I2(n4737), 
            .O(n5405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7194.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7195 (.I0(n5405), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7195.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7196 (.I0(n5405), .I1(n5311), .I2(n5313), .I3(n5406), 
            .O(n17640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7196.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7197 (.I0(\LOAD_DATA[12] ), .I1(\XI[2][12] ), .I2(n4737), 
            .O(n5407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7197.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7198 (.I0(n5407), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7198.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7199 (.I0(n5407), .I1(n5311), .I2(n5313), .I3(n5408), 
            .O(n17639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7199.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7200 (.I0(\LOAD_DATA[13] ), .I1(\XI[2][13] ), .I2(n4737), 
            .O(n5409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7200.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7201 (.I0(n5409), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7201.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7202 (.I0(n5409), .I1(n5311), .I2(n5313), .I3(n5410), 
            .O(n17638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7202.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7203 (.I0(\LOAD_DATA[14] ), .I1(\XI[2][14] ), .I2(n4737), 
            .O(n5411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7203.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7204 (.I0(n5411), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7204.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7205 (.I0(n5411), .I1(n5311), .I2(n5313), .I3(n5412), 
            .O(n17637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7205.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7206 (.I0(\LOAD_DATA[15] ), .I1(\XI[2][15] ), .I2(n4737), 
            .O(n5413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7206.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7207 (.I0(n5413), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7207.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7208 (.I0(n5413), .I1(n5311), .I2(n5313), .I3(n5414), 
            .O(n17636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7208.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7209 (.I0(n4737), .I1(n5330), .O(n5415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7209.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7210 (.I0(\XI[2][16] ), .I1(n5415), .I2(n5334), .I3(n5335), 
            .O(n17635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7210.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7211 (.I0(n4737), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net49837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7211.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7212 (.I0(\XI[2][17] ), .I1(n5415), .I2(n5338), .I3(n5339), 
            .O(n17634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7212.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7213 (.I0(\XI[2][18] ), .I1(n5415), .I2(n5341), .I3(n5342), 
            .O(n17633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7213.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7214 (.I0(\XI[2][19] ), .I1(n5415), .I2(n5344), .I3(n5345), 
            .O(n17632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7214.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7215 (.I0(\XI[2][20] ), .I1(n5415), .I2(n5347), .I3(n5348), 
            .O(n17631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7215.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7216 (.I0(\XI[2][21] ), .I1(n5415), .I2(n5350), .I3(n5351), 
            .O(n17630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7216.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7217 (.I0(\XI[2][22] ), .I1(n5415), .I2(n5353), .I3(n5354), 
            .O(n17629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7217.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7218 (.I0(\XI[2][23] ), .I1(n5415), .I2(n5356), .I3(n5357), 
            .O(n17628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7218.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7219 (.I0(\XI[2][24] ), .I1(n5415), .I2(n5359), .I3(n5360), 
            .O(n17627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7219.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7220 (.I0(\XI[2][25] ), .I1(n5415), .I2(n5362), .I3(n5363), 
            .O(n17626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7220.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7221 (.I0(\XI[2][26] ), .I1(n5415), .I2(n5365), .I3(n5366), 
            .O(n17625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7221.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7222 (.I0(\XI[2][27] ), .I1(n5415), .I2(n5368), .I3(n5369), 
            .O(n17624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7222.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7223 (.I0(\XI[2][28] ), .I1(n5415), .I2(n5371), .I3(n5372), 
            .O(n17623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7223.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7224 (.I0(\XI[2][29] ), .I1(n5415), .I2(n5374), .I3(n5375), 
            .O(n17622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7224.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7225 (.I0(\XI[2][30] ), .I1(n5415), .I2(n5377), .I3(n5378), 
            .O(n17621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7225.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7226 (.I0(\XI[2][31] ), .I1(n5415), .I2(n5380), .I3(n5381), 
            .O(n17620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7226.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7227 (.I0(\LOAD_DATA[8] ), .I1(\XI[3][8] ), .I2(n4739), 
            .O(n5416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7227.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7228 (.I0(n5416), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7228.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7229 (.I0(n5416), .I1(n5311), .I2(n5313), .I3(n5417), 
            .O(n17676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7229.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7230 (.I0(n4739), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net42088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7230.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7231 (.I0(\LOAD_DATA[9] ), .I1(\XI[3][9] ), .I2(n4739), 
            .O(n5418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7231.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7232 (.I0(n5418), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7232.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7233 (.I0(n5418), .I1(n5311), .I2(n5313), .I3(n5419), 
            .O(n17675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7233.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7234 (.I0(\LOAD_DATA[10] ), .I1(\XI[3][10] ), .I2(n4739), 
            .O(n5420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7234.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7235 (.I0(n5420), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7235.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7236 (.I0(n5420), .I1(n5311), .I2(n5313), .I3(n5421), 
            .O(n17674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7236.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7237 (.I0(\LOAD_DATA[11] ), .I1(\XI[3][11] ), .I2(n4739), 
            .O(n5422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7237.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7238 (.I0(n5422), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7238.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7239 (.I0(n5422), .I1(n5311), .I2(n5313), .I3(n5423), 
            .O(n17673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7239.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7240 (.I0(\LOAD_DATA[12] ), .I1(\XI[3][12] ), .I2(n4739), 
            .O(n5424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7240.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7241 (.I0(n5424), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7241.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7242 (.I0(n5424), .I1(n5311), .I2(n5313), .I3(n5425), 
            .O(n17672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7242.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7243 (.I0(\LOAD_DATA[13] ), .I1(\XI[3][13] ), .I2(n4739), 
            .O(n5426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7243.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7244 (.I0(n5426), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7244.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7245 (.I0(n5426), .I1(n5311), .I2(n5313), .I3(n5427), 
            .O(n17671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7245.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7246 (.I0(\LOAD_DATA[14] ), .I1(\XI[3][14] ), .I2(n4739), 
            .O(n5428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7246.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7247 (.I0(n5428), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7247.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7248 (.I0(n5428), .I1(n5311), .I2(n5313), .I3(n5429), 
            .O(n17670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7248.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7249 (.I0(\LOAD_DATA[15] ), .I1(\XI[3][15] ), .I2(n4739), 
            .O(n5430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7249.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7250 (.I0(n5430), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7250.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7251 (.I0(n5430), .I1(n5311), .I2(n5313), .I3(n5431), 
            .O(n17669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7251.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7252 (.I0(n4739), .I1(n5330), .O(n5432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7252.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7253 (.I0(\XI[3][16] ), .I1(n5432), .I2(n5334), .I3(n5335), 
            .O(n17668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7253.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7254 (.I0(n4739), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net49901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7254.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7255 (.I0(\XI[3][17] ), .I1(n5432), .I2(n5338), .I3(n5339), 
            .O(n17667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7255.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7256 (.I0(\XI[3][18] ), .I1(n5432), .I2(n5341), .I3(n5342), 
            .O(n17666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7256.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7257 (.I0(\XI[3][19] ), .I1(n5432), .I2(n5344), .I3(n5345), 
            .O(n17665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7257.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7258 (.I0(\XI[3][20] ), .I1(n5432), .I2(n5347), .I3(n5348), 
            .O(n17664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7258.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7259 (.I0(\XI[3][21] ), .I1(n5432), .I2(n5350), .I3(n5351), 
            .O(n17663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7259.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7260 (.I0(\XI[3][22] ), .I1(n5432), .I2(n5353), .I3(n5354), 
            .O(n17662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7260.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7261 (.I0(\XI[3][23] ), .I1(n5432), .I2(n5356), .I3(n5357), 
            .O(n17661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7261.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7262 (.I0(\XI[3][24] ), .I1(n5432), .I2(n5359), .I3(n5360), 
            .O(n17660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7262.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7263 (.I0(\XI[3][25] ), .I1(n5432), .I2(n5362), .I3(n5363), 
            .O(n17659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7263.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7264 (.I0(\XI[3][26] ), .I1(n5432), .I2(n5365), .I3(n5366), 
            .O(n17658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7264.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7265 (.I0(\XI[3][27] ), .I1(n5432), .I2(n5368), .I3(n5369), 
            .O(n17657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7265.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7266 (.I0(\XI[3][28] ), .I1(n5432), .I2(n5371), .I3(n5372), 
            .O(n17656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7266.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7267 (.I0(\XI[3][29] ), .I1(n5432), .I2(n5374), .I3(n5375), 
            .O(n17655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7267.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7268 (.I0(\XI[3][30] ), .I1(n5432), .I2(n5377), .I3(n5378), 
            .O(n17654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7268.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7269 (.I0(\XI[3][31] ), .I1(n5432), .I2(n5380), .I3(n5381), 
            .O(n17653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7269.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7270 (.I0(\LOAD_DATA[8] ), .I1(\XI[4][8] ), .I2(n4740), 
            .O(n5433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7270.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7271 (.I0(n5433), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7271.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7272 (.I0(n5433), .I1(n5311), .I2(n5313), .I3(n5434), 
            .O(n17709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7272.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7273 (.I0(n4740), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net42280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7273.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7274 (.I0(\LOAD_DATA[9] ), .I1(\XI[4][9] ), .I2(n4740), 
            .O(n5435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7274.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7275 (.I0(n5435), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7275.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7276 (.I0(n5435), .I1(n5311), .I2(n5313), .I3(n5436), 
            .O(n17708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7276.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7277 (.I0(\LOAD_DATA[10] ), .I1(\XI[4][10] ), .I2(n4740), 
            .O(n5437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7277.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7278 (.I0(n5437), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7278.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7279 (.I0(n5437), .I1(n5311), .I2(n5313), .I3(n5438), 
            .O(n17707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7279.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7280 (.I0(\LOAD_DATA[11] ), .I1(\XI[4][11] ), .I2(n4740), 
            .O(n5439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7280.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7281 (.I0(n5439), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7281.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7282 (.I0(n5439), .I1(n5311), .I2(n5313), .I3(n5440), 
            .O(n17706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7282.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7283 (.I0(\LOAD_DATA[12] ), .I1(\XI[4][12] ), .I2(n4740), 
            .O(n5441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7283.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7284 (.I0(n5441), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7284.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7285 (.I0(n5441), .I1(n5311), .I2(n5313), .I3(n5442), 
            .O(n17705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7285.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7286 (.I0(\LOAD_DATA[13] ), .I1(\XI[4][13] ), .I2(n4740), 
            .O(n5443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7286.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7287 (.I0(n5443), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7287.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7288 (.I0(n5443), .I1(n5311), .I2(n5313), .I3(n5444), 
            .O(n17704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7288.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7289 (.I0(\LOAD_DATA[14] ), .I1(\XI[4][14] ), .I2(n4740), 
            .O(n5445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7289.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7290 (.I0(n5445), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7290.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7291 (.I0(n5445), .I1(n5311), .I2(n5313), .I3(n5446), 
            .O(n17703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7291.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7292 (.I0(\LOAD_DATA[15] ), .I1(\XI[4][15] ), .I2(n4740), 
            .O(n5447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7292.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7293 (.I0(n5447), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7293.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7294 (.I0(n5447), .I1(n5311), .I2(n5313), .I3(n5448), 
            .O(n17702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7294.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7295 (.I0(n4740), .I1(n5330), .O(n5449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7295.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7296 (.I0(\XI[4][16] ), .I1(n5449), .I2(n5334), .I3(n5335), 
            .O(n17701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7296.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7297 (.I0(n4740), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net49965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7297.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7298 (.I0(\XI[4][17] ), .I1(n5449), .I2(n5338), .I3(n5339), 
            .O(n17700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7298.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7299 (.I0(\XI[4][18] ), .I1(n5449), .I2(n5341), .I3(n5342), 
            .O(n17699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7299.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7300 (.I0(\XI[4][19] ), .I1(n5449), .I2(n5344), .I3(n5345), 
            .O(n17698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7300.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7301 (.I0(\XI[4][20] ), .I1(n5449), .I2(n5347), .I3(n5348), 
            .O(n17697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7301.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7302 (.I0(\XI[4][21] ), .I1(n5449), .I2(n5350), .I3(n5351), 
            .O(n17696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7302.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7303 (.I0(\XI[4][22] ), .I1(n5449), .I2(n5353), .I3(n5354), 
            .O(n17695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7303.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7304 (.I0(\XI[4][23] ), .I1(n5449), .I2(n5356), .I3(n5357), 
            .O(n17694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7304.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7305 (.I0(\XI[4][24] ), .I1(n5449), .I2(n5359), .I3(n5360), 
            .O(n17693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7305.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7306 (.I0(\XI[4][25] ), .I1(n5449), .I2(n5362), .I3(n5363), 
            .O(n17692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7306.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7307 (.I0(\XI[4][26] ), .I1(n5449), .I2(n5365), .I3(n5366), 
            .O(n17691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7307.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7308 (.I0(\XI[4][27] ), .I1(n5449), .I2(n5368), .I3(n5369), 
            .O(n17690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7308.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7309 (.I0(\XI[4][28] ), .I1(n5449), .I2(n5371), .I3(n5372), 
            .O(n17689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7309.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7310 (.I0(\XI[4][29] ), .I1(n5449), .I2(n5374), .I3(n5375), 
            .O(n17688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7310.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7311 (.I0(\XI[4][30] ), .I1(n5449), .I2(n5377), .I3(n5378), 
            .O(n17687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7311.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7312 (.I0(\XI[4][31] ), .I1(n5449), .I2(n5380), .I3(n5381), 
            .O(n17686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7312.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7313 (.I0(\LOAD_DATA[8] ), .I1(\XI[5][8] ), .I2(n4741), 
            .O(n5450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7313.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7314 (.I0(n5450), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7314.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7315 (.I0(n5450), .I1(n5311), .I2(n5313), .I3(n5451), 
            .O(n17742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7315.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7316 (.I0(n4741), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net42472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7316.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7317 (.I0(\LOAD_DATA[9] ), .I1(\XI[5][9] ), .I2(n4741), 
            .O(n5452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7317.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7318 (.I0(n5452), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7318.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7319 (.I0(n5452), .I1(n5311), .I2(n5313), .I3(n5453), 
            .O(n17741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7319.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7320 (.I0(\LOAD_DATA[10] ), .I1(\XI[5][10] ), .I2(n4741), 
            .O(n5454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7320.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7321 (.I0(n5454), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7321.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7322 (.I0(n5454), .I1(n5311), .I2(n5313), .I3(n5455), 
            .O(n17740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7322.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7323 (.I0(\LOAD_DATA[11] ), .I1(\XI[5][11] ), .I2(n4741), 
            .O(n5456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7323.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7324 (.I0(n5456), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7324.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7325 (.I0(n5456), .I1(n5311), .I2(n5313), .I3(n5457), 
            .O(n17739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7325.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7326 (.I0(\LOAD_DATA[12] ), .I1(\XI[5][12] ), .I2(n4741), 
            .O(n5458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7326.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7327 (.I0(n5458), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7327.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7328 (.I0(n5458), .I1(n5311), .I2(n5313), .I3(n5459), 
            .O(n17738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7328.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7329 (.I0(\LOAD_DATA[13] ), .I1(\XI[5][13] ), .I2(n4741), 
            .O(n5460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7329.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7330 (.I0(n5460), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7330.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7331 (.I0(n5460), .I1(n5311), .I2(n5313), .I3(n5461), 
            .O(n17737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7331.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7332 (.I0(\LOAD_DATA[14] ), .I1(\XI[5][14] ), .I2(n4741), 
            .O(n5462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7332.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7333 (.I0(n5462), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7333.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7334 (.I0(n5462), .I1(n5311), .I2(n5313), .I3(n5463), 
            .O(n17736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7334.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7335 (.I0(\LOAD_DATA[15] ), .I1(\XI[5][15] ), .I2(n4741), 
            .O(n5464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7335.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7336 (.I0(n5464), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7336.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7337 (.I0(n5464), .I1(n5311), .I2(n5313), .I3(n5465), 
            .O(n17735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7337.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7338 (.I0(n4741), .I1(n5330), .O(n5466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7338.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7339 (.I0(\XI[5][16] ), .I1(n5466), .I2(n5334), .I3(n5335), 
            .O(n17734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7339.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7340 (.I0(n4741), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7340.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7341 (.I0(\XI[5][17] ), .I1(n5466), .I2(n5338), .I3(n5339), 
            .O(n17733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7341.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7342 (.I0(\XI[5][18] ), .I1(n5466), .I2(n5341), .I3(n5342), 
            .O(n17732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7342.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7343 (.I0(\XI[5][19] ), .I1(n5466), .I2(n5344), .I3(n5345), 
            .O(n17731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7343.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7344 (.I0(\XI[5][20] ), .I1(n5466), .I2(n5347), .I3(n5348), 
            .O(n17730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7344.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7345 (.I0(\XI[5][21] ), .I1(n5466), .I2(n5350), .I3(n5351), 
            .O(n17729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7345.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7346 (.I0(\XI[5][22] ), .I1(n5466), .I2(n5353), .I3(n5354), 
            .O(n17728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7346.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7347 (.I0(\XI[5][23] ), .I1(n5466), .I2(n5356), .I3(n5357), 
            .O(n17727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7347.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7348 (.I0(\XI[5][24] ), .I1(n5466), .I2(n5359), .I3(n5360), 
            .O(n17726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7348.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7349 (.I0(\XI[5][25] ), .I1(n5466), .I2(n5362), .I3(n5363), 
            .O(n17725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7349.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7350 (.I0(\XI[5][26] ), .I1(n5466), .I2(n5365), .I3(n5366), 
            .O(n17724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7350.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7351 (.I0(\XI[5][27] ), .I1(n5466), .I2(n5368), .I3(n5369), 
            .O(n17723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7351.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7352 (.I0(\XI[5][28] ), .I1(n5466), .I2(n5371), .I3(n5372), 
            .O(n17722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7352.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7353 (.I0(\XI[5][29] ), .I1(n5466), .I2(n5374), .I3(n5375), 
            .O(n17721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7353.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7354 (.I0(\XI[5][30] ), .I1(n5466), .I2(n5377), .I3(n5378), 
            .O(n17720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7354.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7355 (.I0(\XI[5][31] ), .I1(n5466), .I2(n5380), .I3(n5381), 
            .O(n17719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7355.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7356 (.I0(\LOAD_DATA[8] ), .I1(\XI[6][8] ), .I2(n4742), 
            .O(n5467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7356.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7357 (.I0(n5467), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7357.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7358 (.I0(n5467), .I1(n5311), .I2(n5313), .I3(n5468), 
            .O(n17775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7358.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7359 (.I0(n4742), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net42664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7359.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7360 (.I0(\LOAD_DATA[9] ), .I1(\XI[6][9] ), .I2(n4742), 
            .O(n5469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7360.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7361 (.I0(n5469), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7361.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7362 (.I0(n5469), .I1(n5311), .I2(n5313), .I3(n5470), 
            .O(n17774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7362.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7363 (.I0(\LOAD_DATA[10] ), .I1(\XI[6][10] ), .I2(n4742), 
            .O(n5471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7363.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7364 (.I0(n5471), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7364.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7365 (.I0(n5471), .I1(n5311), .I2(n5313), .I3(n5472), 
            .O(n17773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7365.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7366 (.I0(\LOAD_DATA[11] ), .I1(\XI[6][11] ), .I2(n4742), 
            .O(n5473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7366.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7367 (.I0(n5473), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7367.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7368 (.I0(n5473), .I1(n5311), .I2(n5313), .I3(n5474), 
            .O(n17772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7368.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7369 (.I0(\LOAD_DATA[12] ), .I1(\XI[6][12] ), .I2(n4742), 
            .O(n5475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7369.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7370 (.I0(n5475), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7370.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7371 (.I0(n5475), .I1(n5311), .I2(n5313), .I3(n5476), 
            .O(n17771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7371.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7372 (.I0(\LOAD_DATA[13] ), .I1(\XI[6][13] ), .I2(n4742), 
            .O(n5477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7372.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7373 (.I0(n5477), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7373.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7374 (.I0(n5477), .I1(n5311), .I2(n5313), .I3(n5478), 
            .O(n17770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7374.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7375 (.I0(\LOAD_DATA[14] ), .I1(\XI[6][14] ), .I2(n4742), 
            .O(n5479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7375.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7376 (.I0(n5479), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7376.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7377 (.I0(n5479), .I1(n5311), .I2(n5313), .I3(n5480), 
            .O(n17769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7377.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7378 (.I0(\LOAD_DATA[15] ), .I1(\XI[6][15] ), .I2(n4742), 
            .O(n5481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7378.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7379 (.I0(n5481), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7379.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7380 (.I0(n5481), .I1(n5311), .I2(n5313), .I3(n5482), 
            .O(n17768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7380.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7381 (.I0(n4742), .I1(n5330), .O(n5483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7381.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7382 (.I0(\XI[6][16] ), .I1(n5483), .I2(n5334), .I3(n5335), 
            .O(n17767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7382.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7383 (.I0(n4742), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7383.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7384 (.I0(\XI[6][17] ), .I1(n5483), .I2(n5338), .I3(n5339), 
            .O(n17766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7384.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7385 (.I0(\XI[6][18] ), .I1(n5483), .I2(n5341), .I3(n5342), 
            .O(n17765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7385.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7386 (.I0(\XI[6][19] ), .I1(n5483), .I2(n5344), .I3(n5345), 
            .O(n17764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7386.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7387 (.I0(\XI[6][20] ), .I1(n5483), .I2(n5347), .I3(n5348), 
            .O(n17763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7387.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7388 (.I0(\XI[6][21] ), .I1(n5483), .I2(n5350), .I3(n5351), 
            .O(n17762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7388.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7389 (.I0(\XI[6][22] ), .I1(n5483), .I2(n5353), .I3(n5354), 
            .O(n17761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7389.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7390 (.I0(\XI[6][23] ), .I1(n5483), .I2(n5356), .I3(n5357), 
            .O(n17760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7390.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7391 (.I0(\XI[6][24] ), .I1(n5483), .I2(n5359), .I3(n5360), 
            .O(n17759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7391.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7392 (.I0(\XI[6][25] ), .I1(n5483), .I2(n5362), .I3(n5363), 
            .O(n17758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7392.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7393 (.I0(\XI[6][26] ), .I1(n5483), .I2(n5365), .I3(n5366), 
            .O(n17757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7393.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7394 (.I0(\XI[6][27] ), .I1(n5483), .I2(n5368), .I3(n5369), 
            .O(n17756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7394.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7395 (.I0(\XI[6][28] ), .I1(n5483), .I2(n5371), .I3(n5372), 
            .O(n17755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7395.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7396 (.I0(\XI[6][29] ), .I1(n5483), .I2(n5374), .I3(n5375), 
            .O(n17754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7396.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7397 (.I0(\XI[6][30] ), .I1(n5483), .I2(n5377), .I3(n5378), 
            .O(n17753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7397.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7398 (.I0(\XI[6][31] ), .I1(n5483), .I2(n5380), .I3(n5381), 
            .O(n17752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7398.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7399 (.I0(\LOAD_DATA[8] ), .I1(\XI[7][8] ), .I2(n4743), 
            .O(n5484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7399.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7400 (.I0(n5484), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7400.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7401 (.I0(n5484), .I1(n5311), .I2(n5313), .I3(n5485), 
            .O(n17808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7401.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7402 (.I0(n4743), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net42856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7402.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7403 (.I0(\LOAD_DATA[9] ), .I1(\XI[7][9] ), .I2(n4743), 
            .O(n5486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7403.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7404 (.I0(n5486), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7404.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7405 (.I0(n5486), .I1(n5311), .I2(n5313), .I3(n5487), 
            .O(n17807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7405.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7406 (.I0(\LOAD_DATA[10] ), .I1(\XI[7][10] ), .I2(n4743), 
            .O(n5488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7406.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7407 (.I0(n5488), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7407.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7408 (.I0(n5488), .I1(n5311), .I2(n5313), .I3(n5489), 
            .O(n17806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7408.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7409 (.I0(\LOAD_DATA[11] ), .I1(\XI[7][11] ), .I2(n4743), 
            .O(n5490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7409.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7410 (.I0(n5490), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7410.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7411 (.I0(n5490), .I1(n5311), .I2(n5313), .I3(n5491), 
            .O(n17805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7411.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7412 (.I0(\LOAD_DATA[12] ), .I1(\XI[7][12] ), .I2(n4743), 
            .O(n5492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7412.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7413 (.I0(n5492), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7413.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7414 (.I0(n5492), .I1(n5311), .I2(n5313), .I3(n5493), 
            .O(n17804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7414.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7415 (.I0(\LOAD_DATA[13] ), .I1(\XI[7][13] ), .I2(n4743), 
            .O(n5494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7415.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7416 (.I0(n5494), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7416.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7417 (.I0(n5494), .I1(n5311), .I2(n5313), .I3(n5495), 
            .O(n17803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7417.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7418 (.I0(\LOAD_DATA[14] ), .I1(\XI[7][14] ), .I2(n4743), 
            .O(n5496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7418.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7419 (.I0(n5496), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7419.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7420 (.I0(n5496), .I1(n5311), .I2(n5313), .I3(n5497), 
            .O(n17802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7420.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7421 (.I0(\LOAD_DATA[15] ), .I1(\XI[7][15] ), .I2(n4743), 
            .O(n5498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7421.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7422 (.I0(n5498), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7422.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7423 (.I0(n5498), .I1(n5311), .I2(n5313), .I3(n5499), 
            .O(n17801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7423.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7424 (.I0(n4743), .I1(n5330), .O(n5500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7424.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7425 (.I0(\XI[7][16] ), .I1(n5500), .I2(n5334), .I3(n5335), 
            .O(n17800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7425.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7426 (.I0(n4743), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7426.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7427 (.I0(\XI[7][17] ), .I1(n5500), .I2(n5338), .I3(n5339), 
            .O(n17799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7427.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7428 (.I0(\XI[7][18] ), .I1(n5500), .I2(n5341), .I3(n5342), 
            .O(n17798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7428.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7429 (.I0(\XI[7][19] ), .I1(n5500), .I2(n5344), .I3(n5345), 
            .O(n17797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7429.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7430 (.I0(\XI[7][20] ), .I1(n5500), .I2(n5347), .I3(n5348), 
            .O(n17796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7430.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7431 (.I0(\XI[7][21] ), .I1(n5500), .I2(n5350), .I3(n5351), 
            .O(n17795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7431.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7432 (.I0(\XI[7][22] ), .I1(n5500), .I2(n5353), .I3(n5354), 
            .O(n17794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7432.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7433 (.I0(\XI[7][23] ), .I1(n5500), .I2(n5356), .I3(n5357), 
            .O(n17793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7433.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7434 (.I0(\XI[7][24] ), .I1(n5500), .I2(n5359), .I3(n5360), 
            .O(n17792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7434.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7435 (.I0(\XI[7][25] ), .I1(n5500), .I2(n5362), .I3(n5363), 
            .O(n17791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7435.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7436 (.I0(\XI[7][26] ), .I1(n5500), .I2(n5365), .I3(n5366), 
            .O(n17790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7436.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7437 (.I0(\XI[7][27] ), .I1(n5500), .I2(n5368), .I3(n5369), 
            .O(n17789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7437.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7438 (.I0(\XI[7][28] ), .I1(n5500), .I2(n5371), .I3(n5372), 
            .O(n17788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7438.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7439 (.I0(\XI[7][29] ), .I1(n5500), .I2(n5374), .I3(n5375), 
            .O(n17787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7439.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7440 (.I0(\XI[7][30] ), .I1(n5500), .I2(n5377), .I3(n5378), 
            .O(n17786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7440.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7441 (.I0(\XI[7][31] ), .I1(n5500), .I2(n5380), .I3(n5381), 
            .O(n17785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7441.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7442 (.I0(\LOAD_DATA[8] ), .I1(\XI[8][8] ), .I2(n4744), 
            .O(n5501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7442.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7443 (.I0(n5501), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7443.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7444 (.I0(n5501), .I1(n5311), .I2(n5313), .I3(n5502), 
            .O(n17841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7444.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7445 (.I0(n4744), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net43048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7445.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7446 (.I0(\LOAD_DATA[9] ), .I1(\XI[8][9] ), .I2(n4744), 
            .O(n5503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7446.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7447 (.I0(n5503), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7447.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7448 (.I0(n5503), .I1(n5311), .I2(n5313), .I3(n5504), 
            .O(n17840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7448.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7449 (.I0(\LOAD_DATA[10] ), .I1(\XI[8][10] ), .I2(n4744), 
            .O(n5505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7449.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7450 (.I0(n5505), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7450.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7451 (.I0(n5505), .I1(n5311), .I2(n5313), .I3(n5506), 
            .O(n17839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7451.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7452 (.I0(\LOAD_DATA[11] ), .I1(\XI[8][11] ), .I2(n4744), 
            .O(n5507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7452.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7453 (.I0(n5507), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7453.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7454 (.I0(n5507), .I1(n5311), .I2(n5313), .I3(n5508), 
            .O(n17838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7454.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7455 (.I0(\LOAD_DATA[12] ), .I1(\XI[8][12] ), .I2(n4744), 
            .O(n5509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7455.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7456 (.I0(n5509), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7456.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7457 (.I0(n5509), .I1(n5311), .I2(n5313), .I3(n5510), 
            .O(n17837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7457.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7458 (.I0(\LOAD_DATA[13] ), .I1(\XI[8][13] ), .I2(n4744), 
            .O(n5511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7458.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7459 (.I0(n5511), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7459.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7460 (.I0(n5511), .I1(n5311), .I2(n5313), .I3(n5512), 
            .O(n17836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7460.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7461 (.I0(\LOAD_DATA[14] ), .I1(\XI[8][14] ), .I2(n4744), 
            .O(n5513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7461.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7462 (.I0(n5513), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7462.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7463 (.I0(n5513), .I1(n5311), .I2(n5313), .I3(n5514), 
            .O(n17835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7463.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7464 (.I0(\LOAD_DATA[15] ), .I1(\XI[8][15] ), .I2(n4744), 
            .O(n5515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7464.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7465 (.I0(n5515), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7465.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7466 (.I0(n5515), .I1(n5311), .I2(n5313), .I3(n5516), 
            .O(n17834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7466.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7467 (.I0(n4744), .I1(n5330), .O(n5517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7467.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7468 (.I0(\XI[8][16] ), .I1(n5517), .I2(n5334), .I3(n5335), 
            .O(n17833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7468.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7469 (.I0(n4744), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7469.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7470 (.I0(\XI[8][17] ), .I1(n5517), .I2(n5338), .I3(n5339), 
            .O(n17832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7470.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7471 (.I0(\XI[8][18] ), .I1(n5517), .I2(n5341), .I3(n5342), 
            .O(n17831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7471.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7472 (.I0(\XI[8][19] ), .I1(n5517), .I2(n5344), .I3(n5345), 
            .O(n17830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7472.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7473 (.I0(\XI[8][20] ), .I1(n5517), .I2(n5347), .I3(n5348), 
            .O(n17829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7473.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7474 (.I0(\XI[8][21] ), .I1(n5517), .I2(n5350), .I3(n5351), 
            .O(n17828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7474.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7475 (.I0(\XI[8][22] ), .I1(n5517), .I2(n5353), .I3(n5354), 
            .O(n17827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7475.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7476 (.I0(\XI[8][23] ), .I1(n5517), .I2(n5356), .I3(n5357), 
            .O(n17826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7476.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7477 (.I0(\XI[8][24] ), .I1(n5517), .I2(n5359), .I3(n5360), 
            .O(n17825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7477.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7478 (.I0(\XI[8][25] ), .I1(n5517), .I2(n5362), .I3(n5363), 
            .O(n17824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7478.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7479 (.I0(\XI[8][26] ), .I1(n5517), .I2(n5365), .I3(n5366), 
            .O(n17823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7479.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7480 (.I0(\XI[8][27] ), .I1(n5517), .I2(n5368), .I3(n5369), 
            .O(n17822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7480.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7481 (.I0(\XI[8][28] ), .I1(n5517), .I2(n5371), .I3(n5372), 
            .O(n17821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7481.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7482 (.I0(\XI[8][29] ), .I1(n5517), .I2(n5374), .I3(n5375), 
            .O(n17820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7482.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7483 (.I0(\XI[8][30] ), .I1(n5517), .I2(n5377), .I3(n5378), 
            .O(n17819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7483.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7484 (.I0(\XI[8][31] ), .I1(n5517), .I2(n5380), .I3(n5381), 
            .O(n17818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7484.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7485 (.I0(\LOAD_DATA[8] ), .I1(\XI[9][8] ), .I2(n4745), 
            .O(n5518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7485.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7486 (.I0(n5518), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7486.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7487 (.I0(n5518), .I1(n5311), .I2(n5313), .I3(n5519), 
            .O(n17874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7487.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7488 (.I0(n4745), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net43240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7488.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7489 (.I0(\LOAD_DATA[9] ), .I1(\XI[9][9] ), .I2(n4745), 
            .O(n5520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7489.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7490 (.I0(n5520), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7490.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7491 (.I0(n5520), .I1(n5311), .I2(n5313), .I3(n5521), 
            .O(n17873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7491.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7492 (.I0(\LOAD_DATA[10] ), .I1(\XI[9][10] ), .I2(n4745), 
            .O(n5522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7492.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7493 (.I0(n5522), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7493.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7494 (.I0(n5522), .I1(n5311), .I2(n5313), .I3(n5523), 
            .O(n17872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7494.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7495 (.I0(\LOAD_DATA[11] ), .I1(\XI[9][11] ), .I2(n4745), 
            .O(n5524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7495.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7496 (.I0(n5524), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7496.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7497 (.I0(n5524), .I1(n5311), .I2(n5313), .I3(n5525), 
            .O(n17871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7497.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7498 (.I0(\LOAD_DATA[12] ), .I1(\XI[9][12] ), .I2(n4745), 
            .O(n5526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7498.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7499 (.I0(n5526), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7499.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7500 (.I0(n5526), .I1(n5311), .I2(n5313), .I3(n5527), 
            .O(n17870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7500.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7501 (.I0(\LOAD_DATA[13] ), .I1(\XI[9][13] ), .I2(n4745), 
            .O(n5528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7501.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7502 (.I0(n5528), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7502.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7503 (.I0(n5528), .I1(n5311), .I2(n5313), .I3(n5529), 
            .O(n17869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7503.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7504 (.I0(\LOAD_DATA[14] ), .I1(\XI[9][14] ), .I2(n4745), 
            .O(n5530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7504.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7505 (.I0(n5530), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7505.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7506 (.I0(n5530), .I1(n5311), .I2(n5313), .I3(n5531), 
            .O(n17868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7506.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7507 (.I0(\LOAD_DATA[15] ), .I1(\XI[9][15] ), .I2(n4745), 
            .O(n5532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7507.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7508 (.I0(n5532), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7508.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7509 (.I0(n5532), .I1(n5311), .I2(n5313), .I3(n5533), 
            .O(n17867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7509.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7510 (.I0(n4745), .I1(n5330), .O(n5534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7510.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7511 (.I0(\XI[9][16] ), .I1(n5534), .I2(n5334), .I3(n5335), 
            .O(n17866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7511.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7512 (.I0(n4745), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7512.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7513 (.I0(\XI[9][17] ), .I1(n5534), .I2(n5338), .I3(n5339), 
            .O(n17865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7513.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7514 (.I0(\XI[9][18] ), .I1(n5534), .I2(n5341), .I3(n5342), 
            .O(n17864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7514.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7515 (.I0(\XI[9][19] ), .I1(n5534), .I2(n5344), .I3(n5345), 
            .O(n17863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7515.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7516 (.I0(\XI[9][20] ), .I1(n5534), .I2(n5347), .I3(n5348), 
            .O(n17862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7516.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7517 (.I0(\XI[9][21] ), .I1(n5534), .I2(n5350), .I3(n5351), 
            .O(n17861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7517.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7518 (.I0(\XI[9][22] ), .I1(n5534), .I2(n5353), .I3(n5354), 
            .O(n17860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7518.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7519 (.I0(\XI[9][23] ), .I1(n5534), .I2(n5356), .I3(n5357), 
            .O(n17859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7519.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7520 (.I0(\XI[9][24] ), .I1(n5534), .I2(n5359), .I3(n5360), 
            .O(n17858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7520.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7521 (.I0(\XI[9][25] ), .I1(n5534), .I2(n5362), .I3(n5363), 
            .O(n17857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7521.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7522 (.I0(\XI[9][26] ), .I1(n5534), .I2(n5365), .I3(n5366), 
            .O(n17856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7522.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7523 (.I0(\XI[9][27] ), .I1(n5534), .I2(n5368), .I3(n5369), 
            .O(n17855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7523.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7524 (.I0(\XI[9][28] ), .I1(n5534), .I2(n5371), .I3(n5372), 
            .O(n17854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7524.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7525 (.I0(\XI[9][29] ), .I1(n5534), .I2(n5374), .I3(n5375), 
            .O(n17853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7525.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7526 (.I0(\XI[9][30] ), .I1(n5534), .I2(n5377), .I3(n5378), 
            .O(n17852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7526.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7527 (.I0(\XI[9][31] ), .I1(n5534), .I2(n5380), .I3(n5381), 
            .O(n17851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7527.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7528 (.I0(\LOAD_DATA[8] ), .I1(\XI[10][8] ), .I2(n4746), 
            .O(n5535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7528.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7529 (.I0(n5535), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7529.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7530 (.I0(n5535), .I1(n5311), .I2(n5313), .I3(n5536), 
            .O(n17907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7530.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7531 (.I0(n4746), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net43432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7531.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7532 (.I0(\LOAD_DATA[9] ), .I1(\XI[10][9] ), .I2(n4746), 
            .O(n5537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7532.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7533 (.I0(n5537), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7533.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7534 (.I0(n5537), .I1(n5311), .I2(n5313), .I3(n5538), 
            .O(n17906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7534.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7535 (.I0(\LOAD_DATA[10] ), .I1(\XI[10][10] ), .I2(n4746), 
            .O(n5539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7535.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7536 (.I0(n5539), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7536.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7537 (.I0(n5539), .I1(n5311), .I2(n5313), .I3(n5540), 
            .O(n17905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7537.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7538 (.I0(\LOAD_DATA[11] ), .I1(\XI[10][11] ), .I2(n4746), 
            .O(n5541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7538.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7539 (.I0(n5541), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7539.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7540 (.I0(n5541), .I1(n5311), .I2(n5313), .I3(n5542), 
            .O(n17904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7540.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7541 (.I0(\LOAD_DATA[12] ), .I1(\XI[10][12] ), .I2(n4746), 
            .O(n5543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7541.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7542 (.I0(n5543), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7542.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7543 (.I0(n5543), .I1(n5311), .I2(n5313), .I3(n5544), 
            .O(n17903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7543.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7544 (.I0(\LOAD_DATA[13] ), .I1(\XI[10][13] ), .I2(n4746), 
            .O(n5545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7544.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7545 (.I0(n5545), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7545.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7546 (.I0(n5545), .I1(n5311), .I2(n5313), .I3(n5546), 
            .O(n17902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7546.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7547 (.I0(\LOAD_DATA[14] ), .I1(\XI[10][14] ), .I2(n4746), 
            .O(n5547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7547.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7548 (.I0(n5547), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7548.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7549 (.I0(n5547), .I1(n5311), .I2(n5313), .I3(n5548), 
            .O(n17901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7549.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7550 (.I0(\LOAD_DATA[15] ), .I1(\XI[10][15] ), .I2(n4746), 
            .O(n5549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7550.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7551 (.I0(n5549), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7551.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7552 (.I0(n5549), .I1(n5311), .I2(n5313), .I3(n5550), 
            .O(n17900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7552.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7553 (.I0(n4746), .I1(n5330), .O(n5551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7553.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7554 (.I0(\XI[10][16] ), .I1(n5551), .I2(n5334), .I3(n5335), 
            .O(n17899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7554.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7555 (.I0(n4746), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7555.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7556 (.I0(\XI[10][17] ), .I1(n5551), .I2(n5338), .I3(n5339), 
            .O(n17898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7556.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7557 (.I0(\XI[10][18] ), .I1(n5551), .I2(n5341), .I3(n5342), 
            .O(n17897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7557.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7558 (.I0(\XI[10][19] ), .I1(n5551), .I2(n5344), .I3(n5345), 
            .O(n17896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7558.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7559 (.I0(\XI[10][20] ), .I1(n5551), .I2(n5347), .I3(n5348), 
            .O(n17895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7559.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7560 (.I0(\XI[10][21] ), .I1(n5551), .I2(n5350), .I3(n5351), 
            .O(n17894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7560.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7561 (.I0(\XI[10][22] ), .I1(n5551), .I2(n5353), .I3(n5354), 
            .O(n17893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7561.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7562 (.I0(\XI[10][23] ), .I1(n5551), .I2(n5356), .I3(n5357), 
            .O(n17892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7562.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7563 (.I0(\XI[10][24] ), .I1(n5551), .I2(n5359), .I3(n5360), 
            .O(n17891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7563.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7564 (.I0(\XI[10][25] ), .I1(n5551), .I2(n5362), .I3(n5363), 
            .O(n17890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7564.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7565 (.I0(\XI[10][26] ), .I1(n5551), .I2(n5365), .I3(n5366), 
            .O(n17889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7565.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7566 (.I0(\XI[10][27] ), .I1(n5551), .I2(n5368), .I3(n5369), 
            .O(n17888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7566.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7567 (.I0(\XI[10][28] ), .I1(n5551), .I2(n5371), .I3(n5372), 
            .O(n17887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7567.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7568 (.I0(\XI[10][29] ), .I1(n5551), .I2(n5374), .I3(n5375), 
            .O(n17886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7568.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7569 (.I0(\XI[10][30] ), .I1(n5551), .I2(n5377), .I3(n5378), 
            .O(n17885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7569.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7570 (.I0(\XI[10][31] ), .I1(n5551), .I2(n5380), .I3(n5381), 
            .O(n17884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7570.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7571 (.I0(\LOAD_DATA[8] ), .I1(\XI[11][8] ), .I2(n4747), 
            .O(n5552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7571.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7572 (.I0(n5552), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7572.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7573 (.I0(n5552), .I1(n5311), .I2(n5313), .I3(n5553), 
            .O(n17940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7573.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7574 (.I0(n4747), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net43624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7574.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7575 (.I0(\LOAD_DATA[9] ), .I1(\XI[11][9] ), .I2(n4747), 
            .O(n5554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7575.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7576 (.I0(n5554), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7576.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7577 (.I0(n5554), .I1(n5311), .I2(n5313), .I3(n5555), 
            .O(n17939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7577.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7578 (.I0(\LOAD_DATA[10] ), .I1(\XI[11][10] ), .I2(n4747), 
            .O(n5556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7578.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7579 (.I0(n5556), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7579.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7580 (.I0(n5556), .I1(n5311), .I2(n5313), .I3(n5557), 
            .O(n17938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7580.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7581 (.I0(\LOAD_DATA[11] ), .I1(\XI[11][11] ), .I2(n4747), 
            .O(n5558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7581.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7582 (.I0(n5558), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7582.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7583 (.I0(n5558), .I1(n5311), .I2(n5313), .I3(n5559), 
            .O(n17937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7583.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7584 (.I0(\LOAD_DATA[12] ), .I1(\XI[11][12] ), .I2(n4747), 
            .O(n5560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7584.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7585 (.I0(n5560), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7585.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7586 (.I0(n5560), .I1(n5311), .I2(n5313), .I3(n5561), 
            .O(n17936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7586.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7587 (.I0(\LOAD_DATA[13] ), .I1(\XI[11][13] ), .I2(n4747), 
            .O(n5562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7587.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7588 (.I0(n5562), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7588.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7589 (.I0(n5562), .I1(n5311), .I2(n5313), .I3(n5563), 
            .O(n17935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7589.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7590 (.I0(\LOAD_DATA[14] ), .I1(\XI[11][14] ), .I2(n4747), 
            .O(n5564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7590.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7591 (.I0(n5564), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7591.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7592 (.I0(n5564), .I1(n5311), .I2(n5313), .I3(n5565), 
            .O(n17934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7592.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7593 (.I0(\LOAD_DATA[15] ), .I1(\XI[11][15] ), .I2(n4747), 
            .O(n5566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7593.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7594 (.I0(n5566), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7594.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7595 (.I0(n5566), .I1(n5311), .I2(n5313), .I3(n5567), 
            .O(n17933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7595.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7596 (.I0(n4747), .I1(n5330), .O(n5568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7596.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7597 (.I0(\XI[11][16] ), .I1(n5568), .I2(n5334), .I3(n5335), 
            .O(n17932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7597.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7598 (.I0(n4747), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7598.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7599 (.I0(\XI[11][17] ), .I1(n5568), .I2(n5338), .I3(n5339), 
            .O(n17931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7599.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7600 (.I0(\XI[11][18] ), .I1(n5568), .I2(n5341), .I3(n5342), 
            .O(n17930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7600.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7601 (.I0(\XI[11][19] ), .I1(n5568), .I2(n5344), .I3(n5345), 
            .O(n17929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7601.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7602 (.I0(\XI[11][20] ), .I1(n5568), .I2(n5347), .I3(n5348), 
            .O(n17928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7602.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7603 (.I0(\XI[11][21] ), .I1(n5568), .I2(n5350), .I3(n5351), 
            .O(n17927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7603.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7604 (.I0(\XI[11][22] ), .I1(n5568), .I2(n5353), .I3(n5354), 
            .O(n17926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7604.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7605 (.I0(\XI[11][23] ), .I1(n5568), .I2(n5356), .I3(n5357), 
            .O(n17925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7605.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7606 (.I0(\XI[11][24] ), .I1(n5568), .I2(n5359), .I3(n5360), 
            .O(n17924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7606.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7607 (.I0(\XI[11][25] ), .I1(n5568), .I2(n5362), .I3(n5363), 
            .O(n17923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7607.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7608 (.I0(\XI[11][26] ), .I1(n5568), .I2(n5365), .I3(n5366), 
            .O(n17922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7608.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7609 (.I0(\XI[11][27] ), .I1(n5568), .I2(n5368), .I3(n5369), 
            .O(n17921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7609.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7610 (.I0(\XI[11][28] ), .I1(n5568), .I2(n5371), .I3(n5372), 
            .O(n17920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7610.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7611 (.I0(\XI[11][29] ), .I1(n5568), .I2(n5374), .I3(n5375), 
            .O(n17919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7611.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7612 (.I0(\XI[11][30] ), .I1(n5568), .I2(n5377), .I3(n5378), 
            .O(n17918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7612.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7613 (.I0(\XI[11][31] ), .I1(n5568), .I2(n5380), .I3(n5381), 
            .O(n17917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7613.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7614 (.I0(\LOAD_DATA[8] ), .I1(\XI[12][8] ), .I2(n4748), 
            .O(n5569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7614.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7615 (.I0(n5569), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7615.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7616 (.I0(n5569), .I1(n5311), .I2(n5313), .I3(n5570), 
            .O(n17973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7616.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7617 (.I0(n4748), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net43816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7617.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7618 (.I0(\LOAD_DATA[9] ), .I1(\XI[12][9] ), .I2(n4748), 
            .O(n5571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7618.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7619 (.I0(n5571), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7619.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7620 (.I0(n5571), .I1(n5311), .I2(n5313), .I3(n5572), 
            .O(n17972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7620.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7621 (.I0(\LOAD_DATA[10] ), .I1(\XI[12][10] ), .I2(n4748), 
            .O(n5573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7621.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7622 (.I0(n5573), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7622.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7623 (.I0(n5573), .I1(n5311), .I2(n5313), .I3(n5574), 
            .O(n17971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7623.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7624 (.I0(\LOAD_DATA[11] ), .I1(\XI[12][11] ), .I2(n4748), 
            .O(n5575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7624.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7625 (.I0(n5575), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7625.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7626 (.I0(n5575), .I1(n5311), .I2(n5313), .I3(n5576), 
            .O(n17970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7626.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7627 (.I0(\LOAD_DATA[12] ), .I1(\XI[12][12] ), .I2(n4748), 
            .O(n5577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7627.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7628 (.I0(n5577), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7628.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7629 (.I0(n5577), .I1(n5311), .I2(n5313), .I3(n5578), 
            .O(n17969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7629.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7630 (.I0(\LOAD_DATA[13] ), .I1(\XI[12][13] ), .I2(n4748), 
            .O(n5579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7630.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7631 (.I0(n5579), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7631.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7632 (.I0(n5579), .I1(n5311), .I2(n5313), .I3(n5580), 
            .O(n17968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7632.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7633 (.I0(\LOAD_DATA[14] ), .I1(\XI[12][14] ), .I2(n4748), 
            .O(n5581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7633.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7634 (.I0(n5581), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7634.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7635 (.I0(n5581), .I1(n5311), .I2(n5313), .I3(n5582), 
            .O(n17967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7635.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7636 (.I0(\LOAD_DATA[15] ), .I1(\XI[12][15] ), .I2(n4748), 
            .O(n5583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7636.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7637 (.I0(n5583), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7637.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7638 (.I0(n5583), .I1(n5311), .I2(n5313), .I3(n5584), 
            .O(n17966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7638.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7639 (.I0(n4748), .I1(n5330), .O(n5585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7639.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7640 (.I0(\XI[12][16] ), .I1(n5585), .I2(n5334), .I3(n5335), 
            .O(n17965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7640.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7641 (.I0(n4748), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7641.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7642 (.I0(\XI[12][17] ), .I1(n5585), .I2(n5338), .I3(n5339), 
            .O(n17964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7642.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7643 (.I0(\XI[12][18] ), .I1(n5585), .I2(n5341), .I3(n5342), 
            .O(n17963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7643.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7644 (.I0(\XI[12][19] ), .I1(n5585), .I2(n5344), .I3(n5345), 
            .O(n17962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7644.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7645 (.I0(\XI[12][20] ), .I1(n5585), .I2(n5347), .I3(n5348), 
            .O(n17961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7645.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7646 (.I0(\XI[12][21] ), .I1(n5585), .I2(n5350), .I3(n5351), 
            .O(n17960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7646.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7647 (.I0(\XI[12][22] ), .I1(n5585), .I2(n5353), .I3(n5354), 
            .O(n17959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7647.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7648 (.I0(\XI[12][23] ), .I1(n5585), .I2(n5356), .I3(n5357), 
            .O(n17958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7648.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7649 (.I0(\XI[12][24] ), .I1(n5585), .I2(n5359), .I3(n5360), 
            .O(n17957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7649.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7650 (.I0(\XI[12][25] ), .I1(n5585), .I2(n5362), .I3(n5363), 
            .O(n17956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7650.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7651 (.I0(\XI[12][26] ), .I1(n5585), .I2(n5365), .I3(n5366), 
            .O(n17955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7651.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7652 (.I0(\XI[12][27] ), .I1(n5585), .I2(n5368), .I3(n5369), 
            .O(n17954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7652.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7653 (.I0(\XI[12][28] ), .I1(n5585), .I2(n5371), .I3(n5372), 
            .O(n17953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7653.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7654 (.I0(\XI[12][29] ), .I1(n5585), .I2(n5374), .I3(n5375), 
            .O(n17952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7654.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7655 (.I0(\XI[12][30] ), .I1(n5585), .I2(n5377), .I3(n5378), 
            .O(n17951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7655.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7656 (.I0(\XI[12][31] ), .I1(n5585), .I2(n5380), .I3(n5381), 
            .O(n17950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7656.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7657 (.I0(\LOAD_DATA[8] ), .I1(\XI[13][8] ), .I2(n4749), 
            .O(n5586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7657.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7658 (.I0(n5586), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7658.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7659 (.I0(n5586), .I1(n5311), .I2(n5313), .I3(n5587), 
            .O(n18006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7659.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7660 (.I0(n4749), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net44008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7660.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7661 (.I0(\LOAD_DATA[9] ), .I1(\XI[13][9] ), .I2(n4749), 
            .O(n5588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7661.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7662 (.I0(n5588), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7662.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7663 (.I0(n5588), .I1(n5311), .I2(n5313), .I3(n5589), 
            .O(n18005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7663.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7664 (.I0(\LOAD_DATA[10] ), .I1(\XI[13][10] ), .I2(n4749), 
            .O(n5590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7664.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7665 (.I0(n5590), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7665.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7666 (.I0(n5590), .I1(n5311), .I2(n5313), .I3(n5591), 
            .O(n18004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7666.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7667 (.I0(\LOAD_DATA[11] ), .I1(\XI[13][11] ), .I2(n4749), 
            .O(n5592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7667.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7668 (.I0(n5592), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7668.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7669 (.I0(n5592), .I1(n5311), .I2(n5313), .I3(n5593), 
            .O(n18003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7669.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7670 (.I0(\LOAD_DATA[12] ), .I1(\XI[13][12] ), .I2(n4749), 
            .O(n5594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7670.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7671 (.I0(n5594), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7671.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7672 (.I0(n5594), .I1(n5311), .I2(n5313), .I3(n5595), 
            .O(n18002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7672.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7673 (.I0(\LOAD_DATA[13] ), .I1(\XI[13][13] ), .I2(n4749), 
            .O(n5596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7673.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7674 (.I0(n5596), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7674.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7675 (.I0(n5596), .I1(n5311), .I2(n5313), .I3(n5597), 
            .O(n18001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7675.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7676 (.I0(\LOAD_DATA[14] ), .I1(\XI[13][14] ), .I2(n4749), 
            .O(n5598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7676.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7677 (.I0(n5598), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7677.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7678 (.I0(n5598), .I1(n5311), .I2(n5313), .I3(n5599), 
            .O(n18000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7678.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7679 (.I0(\LOAD_DATA[15] ), .I1(\XI[13][15] ), .I2(n4749), 
            .O(n5600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7679.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7680 (.I0(n5600), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7680.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7681 (.I0(n5600), .I1(n5311), .I2(n5313), .I3(n5601), 
            .O(n17999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7681.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7682 (.I0(n4749), .I1(n5330), .O(n5602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7682.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7683 (.I0(\XI[13][16] ), .I1(n5602), .I2(n5334), .I3(n5335), 
            .O(n17998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7683.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7684 (.I0(n4749), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7684.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7685 (.I0(\XI[13][17] ), .I1(n5602), .I2(n5338), .I3(n5339), 
            .O(n17997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7685.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7686 (.I0(\XI[13][18] ), .I1(n5602), .I2(n5341), .I3(n5342), 
            .O(n17996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7686.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7687 (.I0(\XI[13][19] ), .I1(n5602), .I2(n5344), .I3(n5345), 
            .O(n17995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7687.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7688 (.I0(\XI[13][20] ), .I1(n5602), .I2(n5347), .I3(n5348), 
            .O(n17994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7688.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7689 (.I0(\XI[13][21] ), .I1(n5602), .I2(n5350), .I3(n5351), 
            .O(n17993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7689.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7690 (.I0(\XI[13][22] ), .I1(n5602), .I2(n5353), .I3(n5354), 
            .O(n17992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7690.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7691 (.I0(\XI[13][23] ), .I1(n5602), .I2(n5356), .I3(n5357), 
            .O(n17991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7691.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7692 (.I0(\XI[13][24] ), .I1(n5602), .I2(n5359), .I3(n5360), 
            .O(n17990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7692.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7693 (.I0(\XI[13][25] ), .I1(n5602), .I2(n5362), .I3(n5363), 
            .O(n17989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7693.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7694 (.I0(\XI[13][26] ), .I1(n5602), .I2(n5365), .I3(n5366), 
            .O(n17988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7694.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7695 (.I0(\XI[13][27] ), .I1(n5602), .I2(n5368), .I3(n5369), 
            .O(n17987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7695.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7696 (.I0(\XI[13][28] ), .I1(n5602), .I2(n5371), .I3(n5372), 
            .O(n17986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7696.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7697 (.I0(\XI[13][29] ), .I1(n5602), .I2(n5374), .I3(n5375), 
            .O(n17985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7697.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7698 (.I0(\XI[13][30] ), .I1(n5602), .I2(n5377), .I3(n5378), 
            .O(n17984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7698.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7699 (.I0(\XI[13][31] ), .I1(n5602), .I2(n5380), .I3(n5381), 
            .O(n17983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7699.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7700 (.I0(\LOAD_DATA[8] ), .I1(\XI[14][8] ), .I2(n4750), 
            .O(n5603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7700.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7701 (.I0(n5603), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7701.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7702 (.I0(n5603), .I1(n5311), .I2(n5313), .I3(n5604), 
            .O(n18039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7702.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7703 (.I0(n4750), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net44200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7703.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7704 (.I0(\LOAD_DATA[9] ), .I1(\XI[14][9] ), .I2(n4750), 
            .O(n5605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7704.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7705 (.I0(n5605), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7705.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7706 (.I0(n5605), .I1(n5311), .I2(n5313), .I3(n5606), 
            .O(n18038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7706.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7707 (.I0(\LOAD_DATA[10] ), .I1(\XI[14][10] ), .I2(n4750), 
            .O(n5607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7707.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7708 (.I0(n5607), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7708.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7709 (.I0(n5607), .I1(n5311), .I2(n5313), .I3(n5608), 
            .O(n18037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7709.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7710 (.I0(\LOAD_DATA[11] ), .I1(\XI[14][11] ), .I2(n4750), 
            .O(n5609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7710.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7711 (.I0(n5609), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7711.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7712 (.I0(n5609), .I1(n5311), .I2(n5313), .I3(n5610), 
            .O(n18036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7712.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7713 (.I0(\LOAD_DATA[12] ), .I1(\XI[14][12] ), .I2(n4750), 
            .O(n5611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7713.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7714 (.I0(n5611), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7714.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7715 (.I0(n5611), .I1(n5311), .I2(n5313), .I3(n5612), 
            .O(n18035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7715.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7716 (.I0(\LOAD_DATA[13] ), .I1(\XI[14][13] ), .I2(n4750), 
            .O(n5613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7716.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7717 (.I0(n5613), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7717.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7718 (.I0(n5613), .I1(n5311), .I2(n5313), .I3(n5614), 
            .O(n18034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7718.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7719 (.I0(\LOAD_DATA[14] ), .I1(\XI[14][14] ), .I2(n4750), 
            .O(n5615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7719.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7720 (.I0(n5615), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7720.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7721 (.I0(n5615), .I1(n5311), .I2(n5313), .I3(n5616), 
            .O(n18033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7721.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7722 (.I0(\LOAD_DATA[15] ), .I1(\XI[14][15] ), .I2(n4750), 
            .O(n5617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7722.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7723 (.I0(n5617), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7723.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7724 (.I0(n5617), .I1(n5311), .I2(n5313), .I3(n5618), 
            .O(n18032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7724.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7725 (.I0(n4750), .I1(n5330), .O(n5619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7725.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7726 (.I0(\XI[14][16] ), .I1(n5619), .I2(n5334), .I3(n5335), 
            .O(n18031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7726.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7727 (.I0(n4750), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7727.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7728 (.I0(\XI[14][17] ), .I1(n5619), .I2(n5338), .I3(n5339), 
            .O(n18030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7728.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7729 (.I0(\XI[14][18] ), .I1(n5619), .I2(n5341), .I3(n5342), 
            .O(n18029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7729.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7730 (.I0(\XI[14][19] ), .I1(n5619), .I2(n5344), .I3(n5345), 
            .O(n18028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7730.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7731 (.I0(\XI[14][20] ), .I1(n5619), .I2(n5347), .I3(n5348), 
            .O(n18027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7731.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7732 (.I0(\XI[14][21] ), .I1(n5619), .I2(n5350), .I3(n5351), 
            .O(n18026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7732.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7733 (.I0(\XI[14][22] ), .I1(n5619), .I2(n5353), .I3(n5354), 
            .O(n18025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7733.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7734 (.I0(\XI[14][23] ), .I1(n5619), .I2(n5356), .I3(n5357), 
            .O(n18024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7734.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7735 (.I0(\XI[14][24] ), .I1(n5619), .I2(n5359), .I3(n5360), 
            .O(n18023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7735.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7736 (.I0(\XI[14][25] ), .I1(n5619), .I2(n5362), .I3(n5363), 
            .O(n18022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7736.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7737 (.I0(\XI[14][26] ), .I1(n5619), .I2(n5365), .I3(n5366), 
            .O(n18021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7737.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7738 (.I0(\XI[14][27] ), .I1(n5619), .I2(n5368), .I3(n5369), 
            .O(n18020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7738.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7739 (.I0(\XI[14][28] ), .I1(n5619), .I2(n5371), .I3(n5372), 
            .O(n18019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7739.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7740 (.I0(\XI[14][29] ), .I1(n5619), .I2(n5374), .I3(n5375), 
            .O(n18018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7740.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7741 (.I0(\XI[14][30] ), .I1(n5619), .I2(n5377), .I3(n5378), 
            .O(n18017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7741.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7742 (.I0(\XI[14][31] ), .I1(n5619), .I2(n5380), .I3(n5381), 
            .O(n18016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7742.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7743 (.I0(\LOAD_DATA[8] ), .I1(\XI[15][8] ), .I2(n4751), 
            .O(n5620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7743.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7744 (.I0(n5620), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7744.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7745 (.I0(n5620), .I1(n5311), .I2(n5313), .I3(n5621), 
            .O(n18072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7745.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7746 (.I0(n4751), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net44392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7746.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7747 (.I0(\LOAD_DATA[9] ), .I1(\XI[15][9] ), .I2(n4751), 
            .O(n5622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7747.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7748 (.I0(n5622), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7748.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7749 (.I0(n5622), .I1(n5311), .I2(n5313), .I3(n5623), 
            .O(n18071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7749.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7750 (.I0(\LOAD_DATA[10] ), .I1(\XI[15][10] ), .I2(n4751), 
            .O(n5624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7750.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7751 (.I0(n5624), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7751.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7752 (.I0(n5624), .I1(n5311), .I2(n5313), .I3(n5625), 
            .O(n18070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7752.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7753 (.I0(\LOAD_DATA[11] ), .I1(\XI[15][11] ), .I2(n4751), 
            .O(n5626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7753.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7754 (.I0(n5626), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7754.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7755 (.I0(n5626), .I1(n5311), .I2(n5313), .I3(n5627), 
            .O(n18069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7755.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7756 (.I0(\LOAD_DATA[12] ), .I1(\XI[15][12] ), .I2(n4751), 
            .O(n5628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7756.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7757 (.I0(n5628), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7757.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7758 (.I0(n5628), .I1(n5311), .I2(n5313), .I3(n5629), 
            .O(n18068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7758.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7759 (.I0(\LOAD_DATA[13] ), .I1(\XI[15][13] ), .I2(n4751), 
            .O(n5630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7759.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7760 (.I0(n5630), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7760.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7761 (.I0(n5630), .I1(n5311), .I2(n5313), .I3(n5631), 
            .O(n18067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7761.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7762 (.I0(\LOAD_DATA[14] ), .I1(\XI[15][14] ), .I2(n4751), 
            .O(n5632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7762.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7763 (.I0(n5632), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7763.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7764 (.I0(n5632), .I1(n5311), .I2(n5313), .I3(n5633), 
            .O(n18066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7764.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7765 (.I0(\LOAD_DATA[15] ), .I1(\XI[15][15] ), .I2(n4751), 
            .O(n5634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7765.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7766 (.I0(n5634), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7766.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7767 (.I0(n5634), .I1(n5311), .I2(n5313), .I3(n5635), 
            .O(n18065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7767.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7768 (.I0(n4751), .I1(n5330), .O(n5636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7768.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7769 (.I0(\XI[15][16] ), .I1(n5636), .I2(n5334), .I3(n5335), 
            .O(n18064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7769.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7770 (.I0(n4751), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7770.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7771 (.I0(\XI[15][17] ), .I1(n5636), .I2(n5338), .I3(n5339), 
            .O(n18063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7771.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7772 (.I0(\XI[15][18] ), .I1(n5636), .I2(n5341), .I3(n5342), 
            .O(n18062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7772.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7773 (.I0(\XI[15][19] ), .I1(n5636), .I2(n5344), .I3(n5345), 
            .O(n18061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7773.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7774 (.I0(\XI[15][20] ), .I1(n5636), .I2(n5347), .I3(n5348), 
            .O(n18060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7774.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7775 (.I0(\XI[15][21] ), .I1(n5636), .I2(n5350), .I3(n5351), 
            .O(n18059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7775.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7776 (.I0(\XI[15][22] ), .I1(n5636), .I2(n5353), .I3(n5354), 
            .O(n18058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7776.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7777 (.I0(\XI[15][23] ), .I1(n5636), .I2(n5356), .I3(n5357), 
            .O(n18057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7777.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7778 (.I0(\XI[15][24] ), .I1(n5636), .I2(n5359), .I3(n5360), 
            .O(n18056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7778.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7779 (.I0(\XI[15][25] ), .I1(n5636), .I2(n5362), .I3(n5363), 
            .O(n18055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7779.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7780 (.I0(\XI[15][26] ), .I1(n5636), .I2(n5365), .I3(n5366), 
            .O(n18054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7780.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7781 (.I0(\XI[15][27] ), .I1(n5636), .I2(n5368), .I3(n5369), 
            .O(n18053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7781.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7782 (.I0(\XI[15][28] ), .I1(n5636), .I2(n5371), .I3(n5372), 
            .O(n18052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7782.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7783 (.I0(\XI[15][29] ), .I1(n5636), .I2(n5374), .I3(n5375), 
            .O(n18051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7783.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7784 (.I0(\XI[15][30] ), .I1(n5636), .I2(n5377), .I3(n5378), 
            .O(n18050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7784.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7785 (.I0(\XI[15][31] ), .I1(n5636), .I2(n5380), .I3(n5381), 
            .O(n18049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7785.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7786 (.I0(\LOAD_DATA[8] ), .I1(\XI[16][8] ), .I2(n4752), 
            .O(n5637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7786.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7787 (.I0(n5637), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7787.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7788 (.I0(n5637), .I1(n5311), .I2(n5313), .I3(n5638), 
            .O(n18105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7788.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7789 (.I0(n4752), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net44584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7789.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7790 (.I0(\LOAD_DATA[9] ), .I1(\XI[16][9] ), .I2(n4752), 
            .O(n5639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7790.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7791 (.I0(n5639), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7791.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7792 (.I0(n5639), .I1(n5311), .I2(n5313), .I3(n5640), 
            .O(n18104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7792.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7793 (.I0(\LOAD_DATA[10] ), .I1(\XI[16][10] ), .I2(n4752), 
            .O(n5641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7793.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7794 (.I0(n5641), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7794.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7795 (.I0(n5641), .I1(n5311), .I2(n5313), .I3(n5642), 
            .O(n18103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7795.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7796 (.I0(\LOAD_DATA[11] ), .I1(\XI[16][11] ), .I2(n4752), 
            .O(n5643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7796.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7797 (.I0(n5643), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7797.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7798 (.I0(n5643), .I1(n5311), .I2(n5313), .I3(n5644), 
            .O(n18102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7798.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7799 (.I0(\LOAD_DATA[12] ), .I1(\XI[16][12] ), .I2(n4752), 
            .O(n5645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7799.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7800 (.I0(n5645), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7800.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7801 (.I0(n5645), .I1(n5311), .I2(n5313), .I3(n5646), 
            .O(n18101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7801.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7802 (.I0(\LOAD_DATA[13] ), .I1(\XI[16][13] ), .I2(n4752), 
            .O(n5647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7802.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7803 (.I0(n5647), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7803.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7804 (.I0(n5647), .I1(n5311), .I2(n5313), .I3(n5648), 
            .O(n18100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7804.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7805 (.I0(\LOAD_DATA[14] ), .I1(\XI[16][14] ), .I2(n4752), 
            .O(n5649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7805.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7806 (.I0(n5649), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7806.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7807 (.I0(n5649), .I1(n5311), .I2(n5313), .I3(n5650), 
            .O(n18099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7807.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7808 (.I0(\LOAD_DATA[15] ), .I1(\XI[16][15] ), .I2(n4752), 
            .O(n5651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7808.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7809 (.I0(n5651), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7809.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7810 (.I0(n5651), .I1(n5311), .I2(n5313), .I3(n5652), 
            .O(n18098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7810.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7811 (.I0(n4752), .I1(n5330), .O(n5653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7811.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7812 (.I0(\XI[16][16] ), .I1(n5653), .I2(n5334), .I3(n5335), 
            .O(n18097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7812.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7813 (.I0(n4752), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7813.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7814 (.I0(\XI[16][17] ), .I1(n5653), .I2(n5338), .I3(n5339), 
            .O(n18096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7814.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7815 (.I0(\XI[16][18] ), .I1(n5653), .I2(n5341), .I3(n5342), 
            .O(n18095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7815.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7816 (.I0(\XI[16][19] ), .I1(n5653), .I2(n5344), .I3(n5345), 
            .O(n18094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7816.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7817 (.I0(\XI[16][20] ), .I1(n5653), .I2(n5347), .I3(n5348), 
            .O(n18093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7817.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7818 (.I0(\XI[16][21] ), .I1(n5653), .I2(n5350), .I3(n5351), 
            .O(n18092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7818.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7819 (.I0(\XI[16][22] ), .I1(n5653), .I2(n5353), .I3(n5354), 
            .O(n18091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7819.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7820 (.I0(\XI[16][23] ), .I1(n5653), .I2(n5356), .I3(n5357), 
            .O(n18090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7820.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7821 (.I0(\XI[16][24] ), .I1(n5653), .I2(n5359), .I3(n5360), 
            .O(n18089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7821.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7822 (.I0(\XI[16][25] ), .I1(n5653), .I2(n5362), .I3(n5363), 
            .O(n18088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7822.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7823 (.I0(\XI[16][26] ), .I1(n5653), .I2(n5365), .I3(n5366), 
            .O(n18087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7823.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7824 (.I0(\XI[16][27] ), .I1(n5653), .I2(n5368), .I3(n5369), 
            .O(n18086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7824.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7825 (.I0(\XI[16][28] ), .I1(n5653), .I2(n5371), .I3(n5372), 
            .O(n18085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7825.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7826 (.I0(\XI[16][29] ), .I1(n5653), .I2(n5374), .I3(n5375), 
            .O(n18084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7826.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7827 (.I0(\XI[16][30] ), .I1(n5653), .I2(n5377), .I3(n5378), 
            .O(n18083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7827.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7828 (.I0(\XI[16][31] ), .I1(n5653), .I2(n5380), .I3(n5381), 
            .O(n18082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7828.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7829 (.I0(\LOAD_DATA[8] ), .I1(\XI[17][8] ), .I2(n4753), 
            .O(n5654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7829.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7830 (.I0(n5654), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7830.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7831 (.I0(n5654), .I1(n5311), .I2(n5313), .I3(n5655), 
            .O(n18138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7831.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7832 (.I0(n4753), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net44776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7832.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7833 (.I0(\LOAD_DATA[9] ), .I1(\XI[17][9] ), .I2(n4753), 
            .O(n5656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7833.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7834 (.I0(n5656), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7834.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7835 (.I0(n5656), .I1(n5311), .I2(n5313), .I3(n5657), 
            .O(n18137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7835.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7836 (.I0(\LOAD_DATA[10] ), .I1(\XI[17][10] ), .I2(n4753), 
            .O(n5658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7836.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7837 (.I0(n5658), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7837.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7838 (.I0(n5658), .I1(n5311), .I2(n5313), .I3(n5659), 
            .O(n18136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7838.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7839 (.I0(\LOAD_DATA[11] ), .I1(\XI[17][11] ), .I2(n4753), 
            .O(n5660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7839.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7840 (.I0(n5660), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7840.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7841 (.I0(n5660), .I1(n5311), .I2(n5313), .I3(n5661), 
            .O(n18135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7841.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7842 (.I0(\LOAD_DATA[12] ), .I1(\XI[17][12] ), .I2(n4753), 
            .O(n5662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7842.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7843 (.I0(n5662), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7843.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7844 (.I0(n5662), .I1(n5311), .I2(n5313), .I3(n5663), 
            .O(n18134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7844.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7845 (.I0(\LOAD_DATA[13] ), .I1(\XI[17][13] ), .I2(n4753), 
            .O(n5664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7845.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7846 (.I0(n5664), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7846.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7847 (.I0(n5664), .I1(n5311), .I2(n5313), .I3(n5665), 
            .O(n18133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7847.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7848 (.I0(\LOAD_DATA[14] ), .I1(\XI[17][14] ), .I2(n4753), 
            .O(n5666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7848.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7849 (.I0(n5666), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7849.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7850 (.I0(n5666), .I1(n5311), .I2(n5313), .I3(n5667), 
            .O(n18132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7850.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7851 (.I0(\LOAD_DATA[15] ), .I1(\XI[17][15] ), .I2(n4753), 
            .O(n5668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7851.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7852 (.I0(n5668), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7852.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7853 (.I0(n5668), .I1(n5311), .I2(n5313), .I3(n5669), 
            .O(n18131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7853.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7854 (.I0(n4753), .I1(n5330), .O(n5670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7854.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7855 (.I0(\XI[17][16] ), .I1(n5670), .I2(n5334), .I3(n5335), 
            .O(n18130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7855.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7856 (.I0(n4753), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7856.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7857 (.I0(\XI[17][17] ), .I1(n5670), .I2(n5338), .I3(n5339), 
            .O(n18129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7857.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7858 (.I0(\XI[17][18] ), .I1(n5670), .I2(n5341), .I3(n5342), 
            .O(n18128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7858.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7859 (.I0(\XI[17][19] ), .I1(n5670), .I2(n5344), .I3(n5345), 
            .O(n18127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7859.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7860 (.I0(\XI[17][20] ), .I1(n5670), .I2(n5347), .I3(n5348), 
            .O(n18126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7860.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7861 (.I0(\XI[17][21] ), .I1(n5670), .I2(n5350), .I3(n5351), 
            .O(n18125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7861.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7862 (.I0(\XI[17][22] ), .I1(n5670), .I2(n5353), .I3(n5354), 
            .O(n18124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7862.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7863 (.I0(\XI[17][23] ), .I1(n5670), .I2(n5356), .I3(n5357), 
            .O(n18123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7863.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7864 (.I0(\XI[17][24] ), .I1(n5670), .I2(n5359), .I3(n5360), 
            .O(n18122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7864.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7865 (.I0(\XI[17][25] ), .I1(n5670), .I2(n5362), .I3(n5363), 
            .O(n18121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7865.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7866 (.I0(\XI[17][26] ), .I1(n5670), .I2(n5365), .I3(n5366), 
            .O(n18120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7866.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7867 (.I0(\XI[17][27] ), .I1(n5670), .I2(n5368), .I3(n5369), 
            .O(n18119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7867.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7868 (.I0(\XI[17][28] ), .I1(n5670), .I2(n5371), .I3(n5372), 
            .O(n18118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7868.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7869 (.I0(\XI[17][29] ), .I1(n5670), .I2(n5374), .I3(n5375), 
            .O(n18117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7869.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7870 (.I0(\XI[17][30] ), .I1(n5670), .I2(n5377), .I3(n5378), 
            .O(n18116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7870.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7871 (.I0(\XI[17][31] ), .I1(n5670), .I2(n5380), .I3(n5381), 
            .O(n18115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7871.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7872 (.I0(\LOAD_DATA[8] ), .I1(\XI[18][8] ), .I2(n4754), 
            .O(n5671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7872.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7873 (.I0(n5671), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7873.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7874 (.I0(n5671), .I1(n5311), .I2(n5313), .I3(n5672), 
            .O(n18171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7874.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7875 (.I0(n4754), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net44968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7875.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7876 (.I0(\LOAD_DATA[9] ), .I1(\XI[18][9] ), .I2(n4754), 
            .O(n5673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7876.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7877 (.I0(n5673), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7877.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7878 (.I0(n5673), .I1(n5311), .I2(n5313), .I3(n5674), 
            .O(n18170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7878.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7879 (.I0(\LOAD_DATA[10] ), .I1(\XI[18][10] ), .I2(n4754), 
            .O(n5675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7879.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7880 (.I0(n5675), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7880.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7881 (.I0(n5675), .I1(n5311), .I2(n5313), .I3(n5676), 
            .O(n18169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7881.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7882 (.I0(\LOAD_DATA[11] ), .I1(\XI[18][11] ), .I2(n4754), 
            .O(n5677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7882.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7883 (.I0(n5677), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7883.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7884 (.I0(n5677), .I1(n5311), .I2(n5313), .I3(n5678), 
            .O(n18168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7884.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7885 (.I0(\LOAD_DATA[12] ), .I1(\XI[18][12] ), .I2(n4754), 
            .O(n5679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7885.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7886 (.I0(n5679), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7886.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7887 (.I0(n5679), .I1(n5311), .I2(n5313), .I3(n5680), 
            .O(n18167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7887.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7888 (.I0(\LOAD_DATA[13] ), .I1(\XI[18][13] ), .I2(n4754), 
            .O(n5681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7888.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7889 (.I0(n5681), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7889.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7890 (.I0(n5681), .I1(n5311), .I2(n5313), .I3(n5682), 
            .O(n18166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7890.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7891 (.I0(\LOAD_DATA[14] ), .I1(\XI[18][14] ), .I2(n4754), 
            .O(n5683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7891.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7892 (.I0(n5683), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7892.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7893 (.I0(n5683), .I1(n5311), .I2(n5313), .I3(n5684), 
            .O(n18165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7893.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7894 (.I0(\LOAD_DATA[15] ), .I1(\XI[18][15] ), .I2(n4754), 
            .O(n5685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7894.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7895 (.I0(n5685), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7895.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7896 (.I0(n5685), .I1(n5311), .I2(n5313), .I3(n5686), 
            .O(n18164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7896.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7897 (.I0(n4754), .I1(n5330), .O(n5687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7897.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7898 (.I0(\XI[18][16] ), .I1(n5687), .I2(n5334), .I3(n5335), 
            .O(n18163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7898.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7899 (.I0(n4754), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7899.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7900 (.I0(\XI[18][17] ), .I1(n5687), .I2(n5338), .I3(n5339), 
            .O(n18162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7900.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7901 (.I0(\XI[18][18] ), .I1(n5687), .I2(n5341), .I3(n5342), 
            .O(n18161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7901.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7902 (.I0(\XI[18][19] ), .I1(n5687), .I2(n5344), .I3(n5345), 
            .O(n18160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7902.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7903 (.I0(\XI[18][20] ), .I1(n5687), .I2(n5347), .I3(n5348), 
            .O(n18159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7903.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7904 (.I0(\XI[18][21] ), .I1(n5687), .I2(n5350), .I3(n5351), 
            .O(n18158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7904.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7905 (.I0(\XI[18][22] ), .I1(n5687), .I2(n5353), .I3(n5354), 
            .O(n18157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7905.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7906 (.I0(\XI[18][23] ), .I1(n5687), .I2(n5356), .I3(n5357), 
            .O(n18156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7906.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7907 (.I0(\XI[18][24] ), .I1(n5687), .I2(n5359), .I3(n5360), 
            .O(n18155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7907.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7908 (.I0(\XI[18][25] ), .I1(n5687), .I2(n5362), .I3(n5363), 
            .O(n18154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7908.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7909 (.I0(\XI[18][26] ), .I1(n5687), .I2(n5365), .I3(n5366), 
            .O(n18153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7909.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7910 (.I0(\XI[18][27] ), .I1(n5687), .I2(n5368), .I3(n5369), 
            .O(n18152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7910.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7911 (.I0(\XI[18][28] ), .I1(n5687), .I2(n5371), .I3(n5372), 
            .O(n18151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7911.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7912 (.I0(\XI[18][29] ), .I1(n5687), .I2(n5374), .I3(n5375), 
            .O(n18150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7912.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7913 (.I0(\XI[18][30] ), .I1(n5687), .I2(n5377), .I3(n5378), 
            .O(n18149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7913.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7914 (.I0(\XI[18][31] ), .I1(n5687), .I2(n5380), .I3(n5381), 
            .O(n18148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7914.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7915 (.I0(\LOAD_DATA[8] ), .I1(\XI[19][8] ), .I2(n4755), 
            .O(n5688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7915.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7916 (.I0(n5688), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7916.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7917 (.I0(n5688), .I1(n5311), .I2(n5313), .I3(n5689), 
            .O(n18204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7917.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7918 (.I0(n4755), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net45160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7918.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7919 (.I0(\LOAD_DATA[9] ), .I1(\XI[19][9] ), .I2(n4755), 
            .O(n5690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7919.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7920 (.I0(n5690), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7920.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7921 (.I0(n5690), .I1(n5311), .I2(n5313), .I3(n5691), 
            .O(n18203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7921.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7922 (.I0(\LOAD_DATA[10] ), .I1(\XI[19][10] ), .I2(n4755), 
            .O(n5692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7922.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7923 (.I0(n5692), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7923.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7924 (.I0(n5692), .I1(n5311), .I2(n5313), .I3(n5693), 
            .O(n18202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7924.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7925 (.I0(\LOAD_DATA[11] ), .I1(\XI[19][11] ), .I2(n4755), 
            .O(n5694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7925.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7926 (.I0(n5694), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7926.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7927 (.I0(n5694), .I1(n5311), .I2(n5313), .I3(n5695), 
            .O(n18201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7927.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7928 (.I0(\LOAD_DATA[12] ), .I1(\XI[19][12] ), .I2(n4755), 
            .O(n5696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7928.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7929 (.I0(n5696), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7929.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7930 (.I0(n5696), .I1(n5311), .I2(n5313), .I3(n5697), 
            .O(n18200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7930.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7931 (.I0(\LOAD_DATA[13] ), .I1(\XI[19][13] ), .I2(n4755), 
            .O(n5698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7931.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7932 (.I0(n5698), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7932.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7933 (.I0(n5698), .I1(n5311), .I2(n5313), .I3(n5699), 
            .O(n18199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7933.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7934 (.I0(\LOAD_DATA[14] ), .I1(\XI[19][14] ), .I2(n4755), 
            .O(n5700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7934.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7935 (.I0(n5700), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7935.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7936 (.I0(n5700), .I1(n5311), .I2(n5313), .I3(n5701), 
            .O(n18198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7936.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7937 (.I0(\LOAD_DATA[15] ), .I1(\XI[19][15] ), .I2(n4755), 
            .O(n5702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7937.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7938 (.I0(n5702), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7938.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7939 (.I0(n5702), .I1(n5311), .I2(n5313), .I3(n5703), 
            .O(n18197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7939.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7940 (.I0(n4755), .I1(n5330), .O(n5704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7940.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7941 (.I0(\XI[19][16] ), .I1(n5704), .I2(n5334), .I3(n5335), 
            .O(n18196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7941.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7942 (.I0(n4755), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7942.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7943 (.I0(\XI[19][17] ), .I1(n5704), .I2(n5338), .I3(n5339), 
            .O(n18195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7943.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7944 (.I0(\XI[19][18] ), .I1(n5704), .I2(n5341), .I3(n5342), 
            .O(n18194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7944.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7945 (.I0(\XI[19][19] ), .I1(n5704), .I2(n5344), .I3(n5345), 
            .O(n18193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7945.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7946 (.I0(\XI[19][20] ), .I1(n5704), .I2(n5347), .I3(n5348), 
            .O(n18192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7946.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7947 (.I0(\XI[19][21] ), .I1(n5704), .I2(n5350), .I3(n5351), 
            .O(n18191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7947.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7948 (.I0(\XI[19][22] ), .I1(n5704), .I2(n5353), .I3(n5354), 
            .O(n18190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7948.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7949 (.I0(\XI[19][23] ), .I1(n5704), .I2(n5356), .I3(n5357), 
            .O(n18189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7949.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7950 (.I0(\XI[19][24] ), .I1(n5704), .I2(n5359), .I3(n5360), 
            .O(n18188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7950.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7951 (.I0(\XI[19][25] ), .I1(n5704), .I2(n5362), .I3(n5363), 
            .O(n18187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7951.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7952 (.I0(\XI[19][26] ), .I1(n5704), .I2(n5365), .I3(n5366), 
            .O(n18186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7952.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7953 (.I0(\XI[19][27] ), .I1(n5704), .I2(n5368), .I3(n5369), 
            .O(n18185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7953.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7954 (.I0(\XI[19][28] ), .I1(n5704), .I2(n5371), .I3(n5372), 
            .O(n18184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7954.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7955 (.I0(\XI[19][29] ), .I1(n5704), .I2(n5374), .I3(n5375), 
            .O(n18183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7955.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7956 (.I0(\XI[19][30] ), .I1(n5704), .I2(n5377), .I3(n5378), 
            .O(n18182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7956.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7957 (.I0(\XI[19][31] ), .I1(n5704), .I2(n5380), .I3(n5381), 
            .O(n18181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7957.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7958 (.I0(\LOAD_DATA[8] ), .I1(\XI[20][8] ), .I2(n4756), 
            .O(n5705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7958.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7959 (.I0(n5705), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7959.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7960 (.I0(n5705), .I1(n5311), .I2(n5313), .I3(n5706), 
            .O(n18237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7960.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7961 (.I0(n4756), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net45352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7961.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7962 (.I0(\LOAD_DATA[9] ), .I1(\XI[20][9] ), .I2(n4756), 
            .O(n5707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7962.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7963 (.I0(n5707), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7963.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7964 (.I0(n5707), .I1(n5311), .I2(n5313), .I3(n5708), 
            .O(n18236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7964.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7965 (.I0(\LOAD_DATA[10] ), .I1(\XI[20][10] ), .I2(n4756), 
            .O(n5709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7965.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7966 (.I0(n5709), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7966.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7967 (.I0(n5709), .I1(n5311), .I2(n5313), .I3(n5710), 
            .O(n18235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7967.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7968 (.I0(\LOAD_DATA[11] ), .I1(\XI[20][11] ), .I2(n4756), 
            .O(n5711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7968.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7969 (.I0(n5711), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7969.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7970 (.I0(n5711), .I1(n5311), .I2(n5313), .I3(n5712), 
            .O(n18234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7970.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7971 (.I0(\LOAD_DATA[12] ), .I1(\XI[20][12] ), .I2(n4756), 
            .O(n5713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7971.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7972 (.I0(n5713), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7972.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7973 (.I0(n5713), .I1(n5311), .I2(n5313), .I3(n5714), 
            .O(n18233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7973.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7974 (.I0(\LOAD_DATA[13] ), .I1(\XI[20][13] ), .I2(n4756), 
            .O(n5715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7974.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7975 (.I0(n5715), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7975.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7976 (.I0(n5715), .I1(n5311), .I2(n5313), .I3(n5716), 
            .O(n18232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7976.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7977 (.I0(\LOAD_DATA[14] ), .I1(\XI[20][14] ), .I2(n4756), 
            .O(n5717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7977.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7978 (.I0(n5717), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7978.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7979 (.I0(n5717), .I1(n5311), .I2(n5313), .I3(n5718), 
            .O(n18231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7979.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7980 (.I0(\LOAD_DATA[15] ), .I1(\XI[20][15] ), .I2(n4756), 
            .O(n5719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7980.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7981 (.I0(n5719), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__7981.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__7982 (.I0(n5719), .I1(n5311), .I2(n5313), .I3(n5720), 
            .O(n18230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__7982.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__7983 (.I0(n4756), .I1(n5330), .O(n5721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7983.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7984 (.I0(\XI[20][16] ), .I1(n5721), .I2(n5334), .I3(n5335), 
            .O(n18229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7984.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7985 (.I0(n4756), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net50989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__7985.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__7986 (.I0(\XI[20][17] ), .I1(n5721), .I2(n5338), .I3(n5339), 
            .O(n18228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7986.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7987 (.I0(\XI[20][18] ), .I1(n5721), .I2(n5341), .I3(n5342), 
            .O(n18227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7987.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7988 (.I0(\XI[20][19] ), .I1(n5721), .I2(n5344), .I3(n5345), 
            .O(n18226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7988.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7989 (.I0(\XI[20][20] ), .I1(n5721), .I2(n5347), .I3(n5348), 
            .O(n18225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7989.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7990 (.I0(\XI[20][21] ), .I1(n5721), .I2(n5350), .I3(n5351), 
            .O(n18224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7990.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7991 (.I0(\XI[20][22] ), .I1(n5721), .I2(n5353), .I3(n5354), 
            .O(n18223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7991.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7992 (.I0(\XI[20][23] ), .I1(n5721), .I2(n5356), .I3(n5357), 
            .O(n18222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7992.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7993 (.I0(\XI[20][24] ), .I1(n5721), .I2(n5359), .I3(n5360), 
            .O(n18221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7993.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7994 (.I0(\XI[20][25] ), .I1(n5721), .I2(n5362), .I3(n5363), 
            .O(n18220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7994.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7995 (.I0(\XI[20][26] ), .I1(n5721), .I2(n5365), .I3(n5366), 
            .O(n18219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7995.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7996 (.I0(\XI[20][27] ), .I1(n5721), .I2(n5368), .I3(n5369), 
            .O(n18218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7996.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7997 (.I0(\XI[20][28] ), .I1(n5721), .I2(n5371), .I3(n5372), 
            .O(n18217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7997.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7998 (.I0(\XI[20][29] ), .I1(n5721), .I2(n5374), .I3(n5375), 
            .O(n18216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7998.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__7999 (.I0(\XI[20][30] ), .I1(n5721), .I2(n5377), .I3(n5378), 
            .O(n18215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__7999.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8000 (.I0(\XI[20][31] ), .I1(n5721), .I2(n5380), .I3(n5381), 
            .O(n18214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8000.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8001 (.I0(\LOAD_DATA[8] ), .I1(\XI[21][8] ), .I2(n4757), 
            .O(n5722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8001.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8002 (.I0(n5722), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8002.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8003 (.I0(n5722), .I1(n5311), .I2(n5313), .I3(n5723), 
            .O(n18270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8003.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8004 (.I0(n4757), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net45544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8004.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8005 (.I0(\LOAD_DATA[9] ), .I1(\XI[21][9] ), .I2(n4757), 
            .O(n5724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8005.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8006 (.I0(n5724), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8006.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8007 (.I0(n5724), .I1(n5311), .I2(n5313), .I3(n5725), 
            .O(n18269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8007.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8008 (.I0(\LOAD_DATA[10] ), .I1(\XI[21][10] ), .I2(n4757), 
            .O(n5726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8008.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8009 (.I0(n5726), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8009.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8010 (.I0(n5726), .I1(n5311), .I2(n5313), .I3(n5727), 
            .O(n18268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8010.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8011 (.I0(\LOAD_DATA[11] ), .I1(\XI[21][11] ), .I2(n4757), 
            .O(n5728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8011.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8012 (.I0(n5728), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8012.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8013 (.I0(n5728), .I1(n5311), .I2(n5313), .I3(n5729), 
            .O(n18267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8013.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8014 (.I0(\LOAD_DATA[12] ), .I1(\XI[21][12] ), .I2(n4757), 
            .O(n5730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8014.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8015 (.I0(n5730), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8015.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8016 (.I0(n5730), .I1(n5311), .I2(n5313), .I3(n5731), 
            .O(n18266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8016.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8017 (.I0(\LOAD_DATA[13] ), .I1(\XI[21][13] ), .I2(n4757), 
            .O(n5732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8017.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8018 (.I0(n5732), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8018.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8019 (.I0(n5732), .I1(n5311), .I2(n5313), .I3(n5733), 
            .O(n18265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8019.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8020 (.I0(\LOAD_DATA[14] ), .I1(\XI[21][14] ), .I2(n4757), 
            .O(n5734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8020.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8021 (.I0(n5734), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8021.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8022 (.I0(n5734), .I1(n5311), .I2(n5313), .I3(n5735), 
            .O(n18264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8022.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8023 (.I0(\LOAD_DATA[15] ), .I1(\XI[21][15] ), .I2(n4757), 
            .O(n5736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8023.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8024 (.I0(n5736), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8024.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8025 (.I0(n5736), .I1(n5311), .I2(n5313), .I3(n5737), 
            .O(n18263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8025.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8026 (.I0(n4757), .I1(n5330), .O(n5738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8026.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8027 (.I0(\XI[21][16] ), .I1(n5738), .I2(n5334), .I3(n5335), 
            .O(n18262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8027.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8028 (.I0(n4757), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8028.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8029 (.I0(\XI[21][17] ), .I1(n5738), .I2(n5338), .I3(n5339), 
            .O(n18261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8029.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8030 (.I0(\XI[21][18] ), .I1(n5738), .I2(n5341), .I3(n5342), 
            .O(n18260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8030.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8031 (.I0(\XI[21][19] ), .I1(n5738), .I2(n5344), .I3(n5345), 
            .O(n18259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8031.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8032 (.I0(\XI[21][20] ), .I1(n5738), .I2(n5347), .I3(n5348), 
            .O(n18258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8032.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8033 (.I0(\XI[21][21] ), .I1(n5738), .I2(n5350), .I3(n5351), 
            .O(n18257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8033.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8034 (.I0(\XI[21][22] ), .I1(n5738), .I2(n5353), .I3(n5354), 
            .O(n18256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8034.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8035 (.I0(\XI[21][23] ), .I1(n5738), .I2(n5356), .I3(n5357), 
            .O(n18255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8035.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8036 (.I0(\XI[21][24] ), .I1(n5738), .I2(n5359), .I3(n5360), 
            .O(n18254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8036.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8037 (.I0(\XI[21][25] ), .I1(n5738), .I2(n5362), .I3(n5363), 
            .O(n18253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8037.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8038 (.I0(\XI[21][26] ), .I1(n5738), .I2(n5365), .I3(n5366), 
            .O(n18252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8038.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8039 (.I0(\XI[21][27] ), .I1(n5738), .I2(n5368), .I3(n5369), 
            .O(n18251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8039.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8040 (.I0(\XI[21][28] ), .I1(n5738), .I2(n5371), .I3(n5372), 
            .O(n18250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8040.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8041 (.I0(\XI[21][29] ), .I1(n5738), .I2(n5374), .I3(n5375), 
            .O(n18249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8041.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8042 (.I0(\XI[21][30] ), .I1(n5738), .I2(n5377), .I3(n5378), 
            .O(n18248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8042.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8043 (.I0(\XI[21][31] ), .I1(n5738), .I2(n5380), .I3(n5381), 
            .O(n18247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8043.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8044 (.I0(\LOAD_DATA[8] ), .I1(\XI[22][8] ), .I2(n4758), 
            .O(n5739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8044.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8045 (.I0(n5739), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8045.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8046 (.I0(n5739), .I1(n5311), .I2(n5313), .I3(n5740), 
            .O(n18303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8046.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8047 (.I0(n4758), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net45736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8047.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8048 (.I0(\LOAD_DATA[9] ), .I1(\XI[22][9] ), .I2(n4758), 
            .O(n5741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8048.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8049 (.I0(n5741), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8049.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8050 (.I0(n5741), .I1(n5311), .I2(n5313), .I3(n5742), 
            .O(n18302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8050.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8051 (.I0(\LOAD_DATA[10] ), .I1(\XI[22][10] ), .I2(n4758), 
            .O(n5743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8051.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8052 (.I0(n5743), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8052.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8053 (.I0(n5743), .I1(n5311), .I2(n5313), .I3(n5744), 
            .O(n18301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8053.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8054 (.I0(\LOAD_DATA[11] ), .I1(\XI[22][11] ), .I2(n4758), 
            .O(n5745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8054.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8055 (.I0(n5745), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8055.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8056 (.I0(n5745), .I1(n5311), .I2(n5313), .I3(n5746), 
            .O(n18300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8056.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8057 (.I0(\LOAD_DATA[12] ), .I1(\XI[22][12] ), .I2(n4758), 
            .O(n5747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8057.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8058 (.I0(n5747), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8058.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8059 (.I0(n5747), .I1(n5311), .I2(n5313), .I3(n5748), 
            .O(n18299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8059.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8060 (.I0(\LOAD_DATA[13] ), .I1(\XI[22][13] ), .I2(n4758), 
            .O(n5749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8060.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8061 (.I0(n5749), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8061.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8062 (.I0(n5749), .I1(n5311), .I2(n5313), .I3(n5750), 
            .O(n18298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8062.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8063 (.I0(\LOAD_DATA[14] ), .I1(\XI[22][14] ), .I2(n4758), 
            .O(n5751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8063.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8064 (.I0(n5751), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8064.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8065 (.I0(n5751), .I1(n5311), .I2(n5313), .I3(n5752), 
            .O(n18297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8065.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8066 (.I0(\LOAD_DATA[15] ), .I1(\XI[22][15] ), .I2(n4758), 
            .O(n5753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8066.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8067 (.I0(n5753), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8067.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8068 (.I0(n5753), .I1(n5311), .I2(n5313), .I3(n5754), 
            .O(n18296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8068.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8069 (.I0(n4758), .I1(n5330), .O(n5755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8069.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8070 (.I0(\XI[22][16] ), .I1(n5755), .I2(n5334), .I3(n5335), 
            .O(n18295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8070.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8071 (.I0(n4758), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8071.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8072 (.I0(\XI[22][17] ), .I1(n5755), .I2(n5338), .I3(n5339), 
            .O(n18294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8072.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8073 (.I0(\XI[22][18] ), .I1(n5755), .I2(n5341), .I3(n5342), 
            .O(n18293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8073.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8074 (.I0(\XI[22][19] ), .I1(n5755), .I2(n5344), .I3(n5345), 
            .O(n18292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8074.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8075 (.I0(\XI[22][20] ), .I1(n5755), .I2(n5347), .I3(n5348), 
            .O(n18291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8075.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8076 (.I0(\XI[22][21] ), .I1(n5755), .I2(n5350), .I3(n5351), 
            .O(n18290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8076.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8077 (.I0(\XI[22][22] ), .I1(n5755), .I2(n5353), .I3(n5354), 
            .O(n18289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8077.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8078 (.I0(\XI[22][23] ), .I1(n5755), .I2(n5356), .I3(n5357), 
            .O(n18288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8078.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8079 (.I0(\XI[22][24] ), .I1(n5755), .I2(n5359), .I3(n5360), 
            .O(n18287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8079.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8080 (.I0(\XI[22][25] ), .I1(n5755), .I2(n5362), .I3(n5363), 
            .O(n18286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8080.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8081 (.I0(\XI[22][26] ), .I1(n5755), .I2(n5365), .I3(n5366), 
            .O(n18285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8081.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8082 (.I0(\XI[22][27] ), .I1(n5755), .I2(n5368), .I3(n5369), 
            .O(n18284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8082.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8083 (.I0(\XI[22][28] ), .I1(n5755), .I2(n5371), .I3(n5372), 
            .O(n18283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8083.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8084 (.I0(\XI[22][29] ), .I1(n5755), .I2(n5374), .I3(n5375), 
            .O(n18282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8084.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8085 (.I0(\XI[22][30] ), .I1(n5755), .I2(n5377), .I3(n5378), 
            .O(n18281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8085.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8086 (.I0(\XI[22][31] ), .I1(n5755), .I2(n5380), .I3(n5381), 
            .O(n18280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8086.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8087 (.I0(\LOAD_DATA[8] ), .I1(\XI[23][8] ), .I2(n4759), 
            .O(n5756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8087.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8088 (.I0(n5756), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8088.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8089 (.I0(n5756), .I1(n5311), .I2(n5313), .I3(n5757), 
            .O(n18336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8089.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8090 (.I0(n4759), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net45928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8090.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8091 (.I0(\LOAD_DATA[9] ), .I1(\XI[23][9] ), .I2(n4759), 
            .O(n5758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8091.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8092 (.I0(n5758), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8092.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8093 (.I0(n5758), .I1(n5311), .I2(n5313), .I3(n5759), 
            .O(n18335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8093.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8094 (.I0(\LOAD_DATA[10] ), .I1(\XI[23][10] ), .I2(n4759), 
            .O(n5760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8094.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8095 (.I0(n5760), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8095.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8096 (.I0(n5760), .I1(n5311), .I2(n5313), .I3(n5761), 
            .O(n18334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8096.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8097 (.I0(\LOAD_DATA[11] ), .I1(\XI[23][11] ), .I2(n4759), 
            .O(n5762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8097.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8098 (.I0(n5762), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8098.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8099 (.I0(n5762), .I1(n5311), .I2(n5313), .I3(n5763), 
            .O(n18333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8099.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8100 (.I0(\LOAD_DATA[12] ), .I1(\XI[23][12] ), .I2(n4759), 
            .O(n5764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8100.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8101 (.I0(n5764), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8101.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8102 (.I0(n5764), .I1(n5311), .I2(n5313), .I3(n5765), 
            .O(n18332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8102.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8103 (.I0(\LOAD_DATA[13] ), .I1(\XI[23][13] ), .I2(n4759), 
            .O(n5766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8103.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8104 (.I0(n5766), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8104.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8105 (.I0(n5766), .I1(n5311), .I2(n5313), .I3(n5767), 
            .O(n18331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8105.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8106 (.I0(\LOAD_DATA[14] ), .I1(\XI[23][14] ), .I2(n4759), 
            .O(n5768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8106.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8107 (.I0(n5768), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8107.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8108 (.I0(n5768), .I1(n5311), .I2(n5313), .I3(n5769), 
            .O(n18330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8108.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8109 (.I0(\LOAD_DATA[15] ), .I1(\XI[23][15] ), .I2(n4759), 
            .O(n5770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8109.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8110 (.I0(n5770), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8110.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8111 (.I0(n5770), .I1(n5311), .I2(n5313), .I3(n5771), 
            .O(n18329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8111.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8112 (.I0(n4759), .I1(n5330), .O(n5772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8112.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8113 (.I0(\XI[23][16] ), .I1(n5772), .I2(n5334), .I3(n5335), 
            .O(n18328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8113.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8114 (.I0(n4759), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8114.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8115 (.I0(\XI[23][17] ), .I1(n5772), .I2(n5338), .I3(n5339), 
            .O(n18327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8115.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8116 (.I0(\XI[23][18] ), .I1(n5772), .I2(n5341), .I3(n5342), 
            .O(n18326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8116.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8117 (.I0(\XI[23][19] ), .I1(n5772), .I2(n5344), .I3(n5345), 
            .O(n18325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8117.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8118 (.I0(\XI[23][20] ), .I1(n5772), .I2(n5347), .I3(n5348), 
            .O(n18324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8118.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8119 (.I0(\XI[23][21] ), .I1(n5772), .I2(n5350), .I3(n5351), 
            .O(n18323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8119.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8120 (.I0(\XI[23][22] ), .I1(n5772), .I2(n5353), .I3(n5354), 
            .O(n18322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8120.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8121 (.I0(\XI[23][23] ), .I1(n5772), .I2(n5356), .I3(n5357), 
            .O(n18321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8121.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8122 (.I0(\XI[23][24] ), .I1(n5772), .I2(n5359), .I3(n5360), 
            .O(n18320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8122.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8123 (.I0(\XI[23][25] ), .I1(n5772), .I2(n5362), .I3(n5363), 
            .O(n18319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8123.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8124 (.I0(\XI[23][26] ), .I1(n5772), .I2(n5365), .I3(n5366), 
            .O(n18318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8124.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8125 (.I0(\XI[23][27] ), .I1(n5772), .I2(n5368), .I3(n5369), 
            .O(n18317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8125.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8126 (.I0(\XI[23][28] ), .I1(n5772), .I2(n5371), .I3(n5372), 
            .O(n18316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8126.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8127 (.I0(\XI[23][29] ), .I1(n5772), .I2(n5374), .I3(n5375), 
            .O(n18315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8127.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8128 (.I0(\XI[23][30] ), .I1(n5772), .I2(n5377), .I3(n5378), 
            .O(n18314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8128.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8129 (.I0(\XI[23][31] ), .I1(n5772), .I2(n5380), .I3(n5381), 
            .O(n18313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8129.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8130 (.I0(\LOAD_DATA[8] ), .I1(\XI[24][8] ), .I2(n4760), 
            .O(n5773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8130.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8131 (.I0(n5773), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8131.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8132 (.I0(n5773), .I1(n5311), .I2(n5313), .I3(n5774), 
            .O(n18369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8132.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8133 (.I0(n4760), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net46120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8133.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8134 (.I0(\LOAD_DATA[9] ), .I1(\XI[24][9] ), .I2(n4760), 
            .O(n5775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8134.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8135 (.I0(n5775), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8135.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8136 (.I0(n5775), .I1(n5311), .I2(n5313), .I3(n5776), 
            .O(n18368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8136.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8137 (.I0(\LOAD_DATA[10] ), .I1(\XI[24][10] ), .I2(n4760), 
            .O(n5777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8137.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8138 (.I0(n5777), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8138.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8139 (.I0(n5777), .I1(n5311), .I2(n5313), .I3(n5778), 
            .O(n18367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8139.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8140 (.I0(\LOAD_DATA[11] ), .I1(\XI[24][11] ), .I2(n4760), 
            .O(n5779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8140.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8141 (.I0(n5779), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8141.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8142 (.I0(n5779), .I1(n5311), .I2(n5313), .I3(n5780), 
            .O(n18366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8142.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8143 (.I0(\LOAD_DATA[12] ), .I1(\XI[24][12] ), .I2(n4760), 
            .O(n5781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8143.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8144 (.I0(n5781), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8144.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8145 (.I0(n5781), .I1(n5311), .I2(n5313), .I3(n5782), 
            .O(n18365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8145.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8146 (.I0(\LOAD_DATA[13] ), .I1(\XI[24][13] ), .I2(n4760), 
            .O(n5783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8146.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8147 (.I0(n5783), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8147.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8148 (.I0(n5783), .I1(n5311), .I2(n5313), .I3(n5784), 
            .O(n18364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8148.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8149 (.I0(\LOAD_DATA[14] ), .I1(\XI[24][14] ), .I2(n4760), 
            .O(n5785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8149.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8150 (.I0(n5785), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8150.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8151 (.I0(n5785), .I1(n5311), .I2(n5313), .I3(n5786), 
            .O(n18363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8151.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8152 (.I0(\LOAD_DATA[15] ), .I1(\XI[24][15] ), .I2(n4760), 
            .O(n5787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8152.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8153 (.I0(n5787), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8153.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8154 (.I0(n5787), .I1(n5311), .I2(n5313), .I3(n5788), 
            .O(n18362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8154.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8155 (.I0(n4760), .I1(n5330), .O(n5789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8155.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8156 (.I0(\XI[24][16] ), .I1(n5789), .I2(n5334), .I3(n5335), 
            .O(n18361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8156.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8157 (.I0(n4760), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8157.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8158 (.I0(\XI[24][17] ), .I1(n5789), .I2(n5338), .I3(n5339), 
            .O(n18360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8158.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8159 (.I0(\XI[24][18] ), .I1(n5789), .I2(n5341), .I3(n5342), 
            .O(n18359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8159.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8160 (.I0(\XI[24][19] ), .I1(n5789), .I2(n5344), .I3(n5345), 
            .O(n18358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8160.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8161 (.I0(\XI[24][20] ), .I1(n5789), .I2(n5347), .I3(n5348), 
            .O(n18357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8161.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8162 (.I0(\XI[24][21] ), .I1(n5789), .I2(n5350), .I3(n5351), 
            .O(n18356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8162.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8163 (.I0(\XI[24][22] ), .I1(n5789), .I2(n5353), .I3(n5354), 
            .O(n18355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8163.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8164 (.I0(\XI[24][23] ), .I1(n5789), .I2(n5356), .I3(n5357), 
            .O(n18354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8164.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8165 (.I0(\XI[24][24] ), .I1(n5789), .I2(n5359), .I3(n5360), 
            .O(n18353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8165.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8166 (.I0(\XI[24][25] ), .I1(n5789), .I2(n5362), .I3(n5363), 
            .O(n18352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8166.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8167 (.I0(\XI[24][26] ), .I1(n5789), .I2(n5365), .I3(n5366), 
            .O(n18351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8167.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8168 (.I0(\XI[24][27] ), .I1(n5789), .I2(n5368), .I3(n5369), 
            .O(n18350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8168.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8169 (.I0(\XI[24][28] ), .I1(n5789), .I2(n5371), .I3(n5372), 
            .O(n18349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8169.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8170 (.I0(\XI[24][29] ), .I1(n5789), .I2(n5374), .I3(n5375), 
            .O(n18348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8170.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8171 (.I0(\XI[24][30] ), .I1(n5789), .I2(n5377), .I3(n5378), 
            .O(n18347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8171.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8172 (.I0(\XI[24][31] ), .I1(n5789), .I2(n5380), .I3(n5381), 
            .O(n18346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8172.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8173 (.I0(\LOAD_DATA[8] ), .I1(\XI[25][8] ), .I2(n4761), 
            .O(n5790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8173.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8174 (.I0(n5790), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8174.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8175 (.I0(n5790), .I1(n5311), .I2(n5313), .I3(n5791), 
            .O(n18402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8175.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8176 (.I0(n4761), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net46312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8176.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8177 (.I0(\LOAD_DATA[9] ), .I1(\XI[25][9] ), .I2(n4761), 
            .O(n5792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8177.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8178 (.I0(n5792), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8178.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8179 (.I0(n5792), .I1(n5311), .I2(n5313), .I3(n5793), 
            .O(n18401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8179.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8180 (.I0(\LOAD_DATA[10] ), .I1(\XI[25][10] ), .I2(n4761), 
            .O(n5794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8180.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8181 (.I0(n5794), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8181.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8182 (.I0(n5794), .I1(n5311), .I2(n5313), .I3(n5795), 
            .O(n18400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8182.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8183 (.I0(\LOAD_DATA[11] ), .I1(\XI[25][11] ), .I2(n4761), 
            .O(n5796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8183.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8184 (.I0(n5796), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8184.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8185 (.I0(n5796), .I1(n5311), .I2(n5313), .I3(n5797), 
            .O(n18399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8185.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8186 (.I0(\LOAD_DATA[12] ), .I1(\XI[25][12] ), .I2(n4761), 
            .O(n5798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8186.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8187 (.I0(n5798), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8187.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8188 (.I0(n5798), .I1(n5311), .I2(n5313), .I3(n5799), 
            .O(n18398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8188.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8189 (.I0(\LOAD_DATA[13] ), .I1(\XI[25][13] ), .I2(n4761), 
            .O(n5800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8189.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8190 (.I0(n5800), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8190.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8191 (.I0(n5800), .I1(n5311), .I2(n5313), .I3(n5801), 
            .O(n18397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8191.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8192 (.I0(\LOAD_DATA[14] ), .I1(\XI[25][14] ), .I2(n4761), 
            .O(n5802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8192.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8193 (.I0(n5802), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8193.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8194 (.I0(n5802), .I1(n5311), .I2(n5313), .I3(n5803), 
            .O(n18396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8194.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8195 (.I0(\LOAD_DATA[15] ), .I1(\XI[25][15] ), .I2(n4761), 
            .O(n5804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8195.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8196 (.I0(n5804), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8196.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8197 (.I0(n5804), .I1(n5311), .I2(n5313), .I3(n5805), 
            .O(n18395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8197.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8198 (.I0(n4761), .I1(n5330), .O(n5806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8198.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8199 (.I0(\XI[25][16] ), .I1(n5806), .I2(n5334), .I3(n5335), 
            .O(n18394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8199.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8200 (.I0(n4761), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8200.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8201 (.I0(\XI[25][17] ), .I1(n5806), .I2(n5338), .I3(n5339), 
            .O(n18393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8201.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8202 (.I0(\XI[25][18] ), .I1(n5806), .I2(n5341), .I3(n5342), 
            .O(n18392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8202.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8203 (.I0(\XI[25][19] ), .I1(n5806), .I2(n5344), .I3(n5345), 
            .O(n18391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8203.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8204 (.I0(\XI[25][20] ), .I1(n5806), .I2(n5347), .I3(n5348), 
            .O(n18390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8204.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8205 (.I0(\XI[25][21] ), .I1(n5806), .I2(n5350), .I3(n5351), 
            .O(n18389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8205.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8206 (.I0(\XI[25][22] ), .I1(n5806), .I2(n5353), .I3(n5354), 
            .O(n18388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8206.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8207 (.I0(\XI[25][23] ), .I1(n5806), .I2(n5356), .I3(n5357), 
            .O(n18387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8207.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8208 (.I0(\XI[25][24] ), .I1(n5806), .I2(n5359), .I3(n5360), 
            .O(n18386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8208.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8209 (.I0(\XI[25][25] ), .I1(n5806), .I2(n5362), .I3(n5363), 
            .O(n18385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8209.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8210 (.I0(\XI[25][26] ), .I1(n5806), .I2(n5365), .I3(n5366), 
            .O(n18384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8210.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8211 (.I0(\XI[25][27] ), .I1(n5806), .I2(n5368), .I3(n5369), 
            .O(n18383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8211.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8212 (.I0(\XI[25][28] ), .I1(n5806), .I2(n5371), .I3(n5372), 
            .O(n18382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8212.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8213 (.I0(\XI[25][29] ), .I1(n5806), .I2(n5374), .I3(n5375), 
            .O(n18381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8213.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8214 (.I0(\XI[25][30] ), .I1(n5806), .I2(n5377), .I3(n5378), 
            .O(n18380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8214.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8215 (.I0(\XI[25][31] ), .I1(n5806), .I2(n5380), .I3(n5381), 
            .O(n18379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8215.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8216 (.I0(\LOAD_DATA[8] ), .I1(\XI[26][8] ), .I2(n4762), 
            .O(n5807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8216.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8217 (.I0(n5807), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8217.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8218 (.I0(n5807), .I1(n5311), .I2(n5313), .I3(n5808), 
            .O(n18435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8218.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8219 (.I0(n4762), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net46504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8219.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8220 (.I0(\LOAD_DATA[9] ), .I1(\XI[26][9] ), .I2(n4762), 
            .O(n5809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8220.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8221 (.I0(n5809), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8221.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8222 (.I0(n5809), .I1(n5311), .I2(n5313), .I3(n5810), 
            .O(n18434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8222.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8223 (.I0(\LOAD_DATA[10] ), .I1(\XI[26][10] ), .I2(n4762), 
            .O(n5811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8223.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8224 (.I0(n5811), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8224.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8225 (.I0(n5811), .I1(n5311), .I2(n5313), .I3(n5812), 
            .O(n18433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8225.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8226 (.I0(\LOAD_DATA[11] ), .I1(\XI[26][11] ), .I2(n4762), 
            .O(n5813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8226.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8227 (.I0(n5813), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8227.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8228 (.I0(n5813), .I1(n5311), .I2(n5313), .I3(n5814), 
            .O(n18432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8228.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8229 (.I0(\LOAD_DATA[12] ), .I1(\XI[26][12] ), .I2(n4762), 
            .O(n5815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8229.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8230 (.I0(n5815), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8230.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8231 (.I0(n5815), .I1(n5311), .I2(n5313), .I3(n5816), 
            .O(n18431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8231.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8232 (.I0(\LOAD_DATA[13] ), .I1(\XI[26][13] ), .I2(n4762), 
            .O(n5817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8232.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8233 (.I0(n5817), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8233.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8234 (.I0(n5817), .I1(n5311), .I2(n5313), .I3(n5818), 
            .O(n18430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8234.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8235 (.I0(\LOAD_DATA[14] ), .I1(\XI[26][14] ), .I2(n4762), 
            .O(n5819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8235.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8236 (.I0(n5819), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8236.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8237 (.I0(n5819), .I1(n5311), .I2(n5313), .I3(n5820), 
            .O(n18429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8237.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8238 (.I0(\LOAD_DATA[15] ), .I1(\XI[26][15] ), .I2(n4762), 
            .O(n5821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8238.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8239 (.I0(n5821), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8239.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8240 (.I0(n5821), .I1(n5311), .I2(n5313), .I3(n5822), 
            .O(n18428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8240.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8241 (.I0(n4762), .I1(n5330), .O(n5823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8241.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8242 (.I0(\XI[26][16] ), .I1(n5823), .I2(n5334), .I3(n5335), 
            .O(n18427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8242.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8243 (.I0(n4762), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8243.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8244 (.I0(\XI[26][17] ), .I1(n5823), .I2(n5338), .I3(n5339), 
            .O(n18426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8244.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8245 (.I0(\XI[26][18] ), .I1(n5823), .I2(n5341), .I3(n5342), 
            .O(n18425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8245.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8246 (.I0(\XI[26][19] ), .I1(n5823), .I2(n5344), .I3(n5345), 
            .O(n18424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8246.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8247 (.I0(\XI[26][20] ), .I1(n5823), .I2(n5347), .I3(n5348), 
            .O(n18423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8247.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8248 (.I0(\XI[26][21] ), .I1(n5823), .I2(n5350), .I3(n5351), 
            .O(n18422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8248.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8249 (.I0(\XI[26][22] ), .I1(n5823), .I2(n5353), .I3(n5354), 
            .O(n18421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8249.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8250 (.I0(\XI[26][23] ), .I1(n5823), .I2(n5356), .I3(n5357), 
            .O(n18420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8250.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8251 (.I0(\XI[26][24] ), .I1(n5823), .I2(n5359), .I3(n5360), 
            .O(n18419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8251.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8252 (.I0(\XI[26][25] ), .I1(n5823), .I2(n5362), .I3(n5363), 
            .O(n18418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8252.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8253 (.I0(\XI[26][26] ), .I1(n5823), .I2(n5365), .I3(n5366), 
            .O(n18417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8253.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8254 (.I0(\XI[26][27] ), .I1(n5823), .I2(n5368), .I3(n5369), 
            .O(n18416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8254.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8255 (.I0(\XI[26][28] ), .I1(n5823), .I2(n5371), .I3(n5372), 
            .O(n18415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8255.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8256 (.I0(\XI[26][29] ), .I1(n5823), .I2(n5374), .I3(n5375), 
            .O(n18414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8256.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8257 (.I0(\XI[26][30] ), .I1(n5823), .I2(n5377), .I3(n5378), 
            .O(n18413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8257.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8258 (.I0(\XI[26][31] ), .I1(n5823), .I2(n5380), .I3(n5381), 
            .O(n18412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8258.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8259 (.I0(\LOAD_DATA[8] ), .I1(\XI[27][8] ), .I2(n4763), 
            .O(n5824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8259.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8260 (.I0(n5824), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8260.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8261 (.I0(n5824), .I1(n5311), .I2(n5313), .I3(n5825), 
            .O(n18468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8261.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8262 (.I0(n4763), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net46696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8262.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8263 (.I0(\LOAD_DATA[9] ), .I1(\XI[27][9] ), .I2(n4763), 
            .O(n5826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8263.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8264 (.I0(n5826), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8264.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8265 (.I0(n5826), .I1(n5311), .I2(n5313), .I3(n5827), 
            .O(n18467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8265.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8266 (.I0(\LOAD_DATA[10] ), .I1(\XI[27][10] ), .I2(n4763), 
            .O(n5828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8266.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8267 (.I0(n5828), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8267.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8268 (.I0(n5828), .I1(n5311), .I2(n5313), .I3(n5829), 
            .O(n18466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8268.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8269 (.I0(\LOAD_DATA[11] ), .I1(\XI[27][11] ), .I2(n4763), 
            .O(n5830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8269.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8270 (.I0(n5830), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8270.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8271 (.I0(n5830), .I1(n5311), .I2(n5313), .I3(n5831), 
            .O(n18465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8271.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8272 (.I0(\LOAD_DATA[12] ), .I1(\XI[27][12] ), .I2(n4763), 
            .O(n5832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8272.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8273 (.I0(n5832), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8273.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8274 (.I0(n5832), .I1(n5311), .I2(n5313), .I3(n5833), 
            .O(n18464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8274.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8275 (.I0(\LOAD_DATA[13] ), .I1(\XI[27][13] ), .I2(n4763), 
            .O(n5834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8275.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8276 (.I0(n5834), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8276.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8277 (.I0(n5834), .I1(n5311), .I2(n5313), .I3(n5835), 
            .O(n18463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8277.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8278 (.I0(\LOAD_DATA[14] ), .I1(\XI[27][14] ), .I2(n4763), 
            .O(n5836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8278.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8279 (.I0(n5836), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8279.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8280 (.I0(n5836), .I1(n5311), .I2(n5313), .I3(n5837), 
            .O(n18462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8280.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8281 (.I0(\LOAD_DATA[15] ), .I1(\XI[27][15] ), .I2(n4763), 
            .O(n5838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8281.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8282 (.I0(n5838), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8282.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8283 (.I0(n5838), .I1(n5311), .I2(n5313), .I3(n5839), 
            .O(n18461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8283.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8284 (.I0(n4763), .I1(n5330), .O(n5840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8284.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8285 (.I0(\XI[27][16] ), .I1(n5840), .I2(n5334), .I3(n5335), 
            .O(n18460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8285.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8286 (.I0(n4763), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8286.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8287 (.I0(\XI[27][17] ), .I1(n5840), .I2(n5338), .I3(n5339), 
            .O(n18459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8287.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8288 (.I0(\XI[27][18] ), .I1(n5840), .I2(n5341), .I3(n5342), 
            .O(n18458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8288.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8289 (.I0(\XI[27][19] ), .I1(n5840), .I2(n5344), .I3(n5345), 
            .O(n18457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8289.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8290 (.I0(\XI[27][20] ), .I1(n5840), .I2(n5347), .I3(n5348), 
            .O(n18456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8290.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8291 (.I0(\XI[27][21] ), .I1(n5840), .I2(n5350), .I3(n5351), 
            .O(n18455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8291.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8292 (.I0(\XI[27][22] ), .I1(n5840), .I2(n5353), .I3(n5354), 
            .O(n18454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8292.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8293 (.I0(\XI[27][23] ), .I1(n5840), .I2(n5356), .I3(n5357), 
            .O(n18453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8293.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8294 (.I0(\XI[27][24] ), .I1(n5840), .I2(n5359), .I3(n5360), 
            .O(n18452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8294.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8295 (.I0(\XI[27][25] ), .I1(n5840), .I2(n5362), .I3(n5363), 
            .O(n18451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8295.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8296 (.I0(\XI[27][26] ), .I1(n5840), .I2(n5365), .I3(n5366), 
            .O(n18450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8296.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8297 (.I0(\XI[27][27] ), .I1(n5840), .I2(n5368), .I3(n5369), 
            .O(n18449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8297.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8298 (.I0(\XI[27][28] ), .I1(n5840), .I2(n5371), .I3(n5372), 
            .O(n18448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8298.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8299 (.I0(\XI[27][29] ), .I1(n5840), .I2(n5374), .I3(n5375), 
            .O(n18447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8299.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8300 (.I0(\XI[27][30] ), .I1(n5840), .I2(n5377), .I3(n5378), 
            .O(n18446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8300.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8301 (.I0(\XI[27][31] ), .I1(n5840), .I2(n5380), .I3(n5381), 
            .O(n18445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8301.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8302 (.I0(\LOAD_DATA[8] ), .I1(\XI[28][8] ), .I2(n4764), 
            .O(n5841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8302.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8303 (.I0(n5841), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8303.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8304 (.I0(n5841), .I1(n5311), .I2(n5313), .I3(n5842), 
            .O(n18501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8304.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8305 (.I0(n4764), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net46888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8305.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8306 (.I0(\LOAD_DATA[9] ), .I1(\XI[28][9] ), .I2(n4764), 
            .O(n5843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8306.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8307 (.I0(n5843), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8307.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8308 (.I0(n5843), .I1(n5311), .I2(n5313), .I3(n5844), 
            .O(n18500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8308.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8309 (.I0(\LOAD_DATA[10] ), .I1(\XI[28][10] ), .I2(n4764), 
            .O(n5845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8309.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8310 (.I0(n5845), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8310.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8311 (.I0(n5845), .I1(n5311), .I2(n5313), .I3(n5846), 
            .O(n18499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8311.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8312 (.I0(\LOAD_DATA[11] ), .I1(\XI[28][11] ), .I2(n4764), 
            .O(n5847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8312.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8313 (.I0(n5847), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8313.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8314 (.I0(n5847), .I1(n5311), .I2(n5313), .I3(n5848), 
            .O(n18498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8314.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8315 (.I0(\LOAD_DATA[12] ), .I1(\XI[28][12] ), .I2(n4764), 
            .O(n5849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8315.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8316 (.I0(n5849), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8316.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8317 (.I0(n5849), .I1(n5311), .I2(n5313), .I3(n5850), 
            .O(n18497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8317.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8318 (.I0(\LOAD_DATA[13] ), .I1(\XI[28][13] ), .I2(n4764), 
            .O(n5851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8318.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8319 (.I0(n5851), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8319.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8320 (.I0(n5851), .I1(n5311), .I2(n5313), .I3(n5852), 
            .O(n18496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8320.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8321 (.I0(\LOAD_DATA[14] ), .I1(\XI[28][14] ), .I2(n4764), 
            .O(n5853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8321.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8322 (.I0(n5853), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8322.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8323 (.I0(n5853), .I1(n5311), .I2(n5313), .I3(n5854), 
            .O(n18495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8323.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8324 (.I0(\LOAD_DATA[15] ), .I1(\XI[28][15] ), .I2(n4764), 
            .O(n5855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8324.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8325 (.I0(n5855), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8325.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8326 (.I0(n5855), .I1(n5311), .I2(n5313), .I3(n5856), 
            .O(n18494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8326.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8327 (.I0(n4764), .I1(n5330), .O(n5857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8327.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8328 (.I0(\XI[28][16] ), .I1(n5857), .I2(n5334), .I3(n5335), 
            .O(n18493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8328.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8329 (.I0(n4764), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8329.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8330 (.I0(\XI[28][17] ), .I1(n5857), .I2(n5338), .I3(n5339), 
            .O(n18492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8330.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8331 (.I0(\XI[28][18] ), .I1(n5857), .I2(n5341), .I3(n5342), 
            .O(n18491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8331.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8332 (.I0(\XI[28][19] ), .I1(n5857), .I2(n5344), .I3(n5345), 
            .O(n18490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8332.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8333 (.I0(\XI[28][20] ), .I1(n5857), .I2(n5347), .I3(n5348), 
            .O(n18489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8333.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8334 (.I0(\XI[28][21] ), .I1(n5857), .I2(n5350), .I3(n5351), 
            .O(n18488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8334.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8335 (.I0(\XI[28][22] ), .I1(n5857), .I2(n5353), .I3(n5354), 
            .O(n18487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8335.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8336 (.I0(\XI[28][23] ), .I1(n5857), .I2(n5356), .I3(n5357), 
            .O(n18486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8336.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8337 (.I0(\XI[28][24] ), .I1(n5857), .I2(n5359), .I3(n5360), 
            .O(n18485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8337.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8338 (.I0(\XI[28][25] ), .I1(n5857), .I2(n5362), .I3(n5363), 
            .O(n18484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8338.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8339 (.I0(\XI[28][26] ), .I1(n5857), .I2(n5365), .I3(n5366), 
            .O(n18483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8339.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8340 (.I0(\XI[28][27] ), .I1(n5857), .I2(n5368), .I3(n5369), 
            .O(n18482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8340.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8341 (.I0(\XI[28][28] ), .I1(n5857), .I2(n5371), .I3(n5372), 
            .O(n18481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8341.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8342 (.I0(\XI[28][29] ), .I1(n5857), .I2(n5374), .I3(n5375), 
            .O(n18480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8342.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8343 (.I0(\XI[28][30] ), .I1(n5857), .I2(n5377), .I3(n5378), 
            .O(n18479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8343.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8344 (.I0(\XI[28][31] ), .I1(n5857), .I2(n5380), .I3(n5381), 
            .O(n18478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8344.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8345 (.I0(\LOAD_DATA[8] ), .I1(\XI[29][8] ), .I2(n4765), 
            .O(n5858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8345.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8346 (.I0(n5858), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8346.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8347 (.I0(n5858), .I1(n5311), .I2(n5313), .I3(n5859), 
            .O(n18534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8347.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8348 (.I0(n4765), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net47080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8348.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8349 (.I0(\LOAD_DATA[9] ), .I1(\XI[29][9] ), .I2(n4765), 
            .O(n5860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8349.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8350 (.I0(n5860), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8350.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8351 (.I0(n5860), .I1(n5311), .I2(n5313), .I3(n5861), 
            .O(n18533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8351.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8352 (.I0(\LOAD_DATA[10] ), .I1(\XI[29][10] ), .I2(n4765), 
            .O(n5862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8352.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8353 (.I0(n5862), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8353.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8354 (.I0(n5862), .I1(n5311), .I2(n5313), .I3(n5863), 
            .O(n18532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8354.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8355 (.I0(\LOAD_DATA[11] ), .I1(\XI[29][11] ), .I2(n4765), 
            .O(n5864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8355.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8356 (.I0(n5864), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8356.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8357 (.I0(n5864), .I1(n5311), .I2(n5313), .I3(n5865), 
            .O(n18531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8357.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8358 (.I0(\LOAD_DATA[12] ), .I1(\XI[29][12] ), .I2(n4765), 
            .O(n5866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8358.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8359 (.I0(n5866), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8359.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8360 (.I0(n5866), .I1(n5311), .I2(n5313), .I3(n5867), 
            .O(n18530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8360.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8361 (.I0(\LOAD_DATA[13] ), .I1(\XI[29][13] ), .I2(n4765), 
            .O(n5868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8361.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8362 (.I0(n5868), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8362.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8363 (.I0(n5868), .I1(n5311), .I2(n5313), .I3(n5869), 
            .O(n18529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8363.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8364 (.I0(\LOAD_DATA[14] ), .I1(\XI[29][14] ), .I2(n4765), 
            .O(n5870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8364.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8365 (.I0(n5870), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8365.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8366 (.I0(n5870), .I1(n5311), .I2(n5313), .I3(n5871), 
            .O(n18528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8366.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8367 (.I0(\LOAD_DATA[15] ), .I1(\XI[29][15] ), .I2(n4765), 
            .O(n5872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8367.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8368 (.I0(n5872), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8368.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8369 (.I0(n5872), .I1(n5311), .I2(n5313), .I3(n5873), 
            .O(n18527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8369.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8370 (.I0(n4765), .I1(n5330), .O(n5874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8370.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8371 (.I0(\XI[29][16] ), .I1(n5874), .I2(n5334), .I3(n5335), 
            .O(n18526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8371.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8372 (.I0(n4765), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8372.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8373 (.I0(\XI[29][17] ), .I1(n5874), .I2(n5338), .I3(n5339), 
            .O(n18525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8373.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8374 (.I0(\XI[29][18] ), .I1(n5874), .I2(n5341), .I3(n5342), 
            .O(n18524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8374.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8375 (.I0(\XI[29][19] ), .I1(n5874), .I2(n5344), .I3(n5345), 
            .O(n18523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8375.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8376 (.I0(\XI[29][20] ), .I1(n5874), .I2(n5347), .I3(n5348), 
            .O(n18522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8376.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8377 (.I0(\XI[29][21] ), .I1(n5874), .I2(n5350), .I3(n5351), 
            .O(n18521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8377.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8378 (.I0(\XI[29][22] ), .I1(n5874), .I2(n5353), .I3(n5354), 
            .O(n18520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8378.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8379 (.I0(\XI[29][23] ), .I1(n5874), .I2(n5356), .I3(n5357), 
            .O(n18519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8379.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8380 (.I0(\XI[29][24] ), .I1(n5874), .I2(n5359), .I3(n5360), 
            .O(n18518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8380.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8381 (.I0(\XI[29][25] ), .I1(n5874), .I2(n5362), .I3(n5363), 
            .O(n18517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8381.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8382 (.I0(\XI[29][26] ), .I1(n5874), .I2(n5365), .I3(n5366), 
            .O(n18516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8382.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8383 (.I0(\XI[29][27] ), .I1(n5874), .I2(n5368), .I3(n5369), 
            .O(n18515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8383.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8384 (.I0(\XI[29][28] ), .I1(n5874), .I2(n5371), .I3(n5372), 
            .O(n18514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8384.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8385 (.I0(\XI[29][29] ), .I1(n5874), .I2(n5374), .I3(n5375), 
            .O(n18513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8385.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8386 (.I0(\XI[29][30] ), .I1(n5874), .I2(n5377), .I3(n5378), 
            .O(n18512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8386.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8387 (.I0(\XI[29][31] ), .I1(n5874), .I2(n5380), .I3(n5381), 
            .O(n18511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8387.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8388 (.I0(\LOAD_DATA[8] ), .I1(\XI[30][8] ), .I2(n4766), 
            .O(n5875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8388.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8389 (.I0(n5875), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8389.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8390 (.I0(n5875), .I1(n5311), .I2(n5313), .I3(n5876), 
            .O(n18567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8390.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8391 (.I0(n4766), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net47272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8391.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8392 (.I0(\LOAD_DATA[9] ), .I1(\XI[30][9] ), .I2(n4766), 
            .O(n5877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8392.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8393 (.I0(n5877), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8393.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8394 (.I0(n5877), .I1(n5311), .I2(n5313), .I3(n5878), 
            .O(n18566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8394.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8395 (.I0(\LOAD_DATA[10] ), .I1(\XI[30][10] ), .I2(n4766), 
            .O(n5879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8395.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8396 (.I0(n5879), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8396.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8397 (.I0(n5879), .I1(n5311), .I2(n5313), .I3(n5880), 
            .O(n18565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8397.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8398 (.I0(\LOAD_DATA[11] ), .I1(\XI[30][11] ), .I2(n4766), 
            .O(n5881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8398.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8399 (.I0(n5881), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8399.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8400 (.I0(n5881), .I1(n5311), .I2(n5313), .I3(n5882), 
            .O(n18564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8400.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8401 (.I0(\LOAD_DATA[12] ), .I1(\XI[30][12] ), .I2(n4766), 
            .O(n5883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8401.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8402 (.I0(n5883), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8402.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8403 (.I0(n5883), .I1(n5311), .I2(n5313), .I3(n5884), 
            .O(n18563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8403.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8404 (.I0(\LOAD_DATA[13] ), .I1(\XI[30][13] ), .I2(n4766), 
            .O(n5885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8404.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8405 (.I0(n5885), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8405.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8406 (.I0(n5885), .I1(n5311), .I2(n5313), .I3(n5886), 
            .O(n18562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8406.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8407 (.I0(\LOAD_DATA[14] ), .I1(\XI[30][14] ), .I2(n4766), 
            .O(n5887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8407.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8408 (.I0(n5887), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8408.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8409 (.I0(n5887), .I1(n5311), .I2(n5313), .I3(n5888), 
            .O(n18561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8409.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8410 (.I0(\LOAD_DATA[15] ), .I1(\XI[30][15] ), .I2(n4766), 
            .O(n5889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8410.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8411 (.I0(n5889), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8411.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8412 (.I0(n5889), .I1(n5311), .I2(n5313), .I3(n5890), 
            .O(n18560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8412.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8413 (.I0(n4766), .I1(n5330), .O(n5891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8413.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8414 (.I0(\XI[30][16] ), .I1(n5891), .I2(n5334), .I3(n5335), 
            .O(n18559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8414.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8415 (.I0(n4766), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8415.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8416 (.I0(\XI[30][17] ), .I1(n5891), .I2(n5338), .I3(n5339), 
            .O(n18558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8416.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8417 (.I0(\XI[30][18] ), .I1(n5891), .I2(n5341), .I3(n5342), 
            .O(n18557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8417.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8418 (.I0(\XI[30][19] ), .I1(n5891), .I2(n5344), .I3(n5345), 
            .O(n18556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8418.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8419 (.I0(\XI[30][20] ), .I1(n5891), .I2(n5347), .I3(n5348), 
            .O(n18555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8419.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8420 (.I0(\XI[30][21] ), .I1(n5891), .I2(n5350), .I3(n5351), 
            .O(n18554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8420.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8421 (.I0(\XI[30][22] ), .I1(n5891), .I2(n5353), .I3(n5354), 
            .O(n18553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8421.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8422 (.I0(\XI[30][23] ), .I1(n5891), .I2(n5356), .I3(n5357), 
            .O(n18552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8422.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8423 (.I0(\XI[30][24] ), .I1(n5891), .I2(n5359), .I3(n5360), 
            .O(n18551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8423.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8424 (.I0(\XI[30][25] ), .I1(n5891), .I2(n5362), .I3(n5363), 
            .O(n18550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8424.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8425 (.I0(\XI[30][26] ), .I1(n5891), .I2(n5365), .I3(n5366), 
            .O(n18549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8425.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8426 (.I0(\XI[30][27] ), .I1(n5891), .I2(n5368), .I3(n5369), 
            .O(n18548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8426.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8427 (.I0(\XI[30][28] ), .I1(n5891), .I2(n5371), .I3(n5372), 
            .O(n18547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8427.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8428 (.I0(\XI[30][29] ), .I1(n5891), .I2(n5374), .I3(n5375), 
            .O(n18546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8428.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8429 (.I0(\XI[30][30] ), .I1(n5891), .I2(n5377), .I3(n5378), 
            .O(n18545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8429.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8430 (.I0(\XI[30][31] ), .I1(n5891), .I2(n5380), .I3(n5381), 
            .O(n18544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8430.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8431 (.I0(\LOAD_DATA[8] ), .I1(\XI[31][8] ), .I2(n4767), 
            .O(n5892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8431.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8432 (.I0(n5892), .I1(n1607), .I2(n5312), .I3(n5310), 
            .O(n5893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8432.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8433 (.I0(n5892), .I1(n5311), .I2(n5313), .I3(n5893), 
            .O(n18600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8433.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8434 (.I0(n4767), .I1(n5315), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net47464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8434.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8435 (.I0(\LOAD_DATA[9] ), .I1(\XI[31][9] ), .I2(n4767), 
            .O(n5894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8435.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8436 (.I0(n5894), .I1(n1606), .I2(n5312), .I3(n5310), 
            .O(n5895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8436.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8437 (.I0(n5894), .I1(n5311), .I2(n5313), .I3(n5895), 
            .O(n18599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8437.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8438 (.I0(\LOAD_DATA[10] ), .I1(\XI[31][10] ), .I2(n4767), 
            .O(n5896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8438.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8439 (.I0(n5896), .I1(n1605), .I2(n5312), .I3(n5310), 
            .O(n5897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8439.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8440 (.I0(n5896), .I1(n5311), .I2(n5313), .I3(n5897), 
            .O(n18598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8440.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8441 (.I0(\LOAD_DATA[11] ), .I1(\XI[31][11] ), .I2(n4767), 
            .O(n5898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8441.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8442 (.I0(n5898), .I1(n1604), .I2(n5312), .I3(n5310), 
            .O(n5899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8442.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8443 (.I0(n5898), .I1(n5311), .I2(n5313), .I3(n5899), 
            .O(n18597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8443.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8444 (.I0(\LOAD_DATA[12] ), .I1(\XI[31][12] ), .I2(n4767), 
            .O(n5900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8444.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8445 (.I0(n5900), .I1(n1603_2), .I2(n5312), .I3(n5310), 
            .O(n5901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8445.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8446 (.I0(n5900), .I1(n5311), .I2(n5313), .I3(n5901), 
            .O(n18596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8446.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8447 (.I0(\LOAD_DATA[13] ), .I1(\XI[31][13] ), .I2(n4767), 
            .O(n5902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8447.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8448 (.I0(n5902), .I1(n1602_2), .I2(n5312), .I3(n5310), 
            .O(n5903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8448.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8449 (.I0(n5902), .I1(n5311), .I2(n5313), .I3(n5903), 
            .O(n18595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8449.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8450 (.I0(\LOAD_DATA[14] ), .I1(\XI[31][14] ), .I2(n4767), 
            .O(n5904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8450.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8451 (.I0(n5904), .I1(n1601_2), .I2(n5312), .I3(n5310), 
            .O(n5905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8451.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8452 (.I0(n5904), .I1(n5311), .I2(n5313), .I3(n5905), 
            .O(n18594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8452.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8453 (.I0(\LOAD_DATA[15] ), .I1(\XI[31][15] ), .I2(n4767), 
            .O(n5906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8453.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8454 (.I0(n5906), .I1(n1600_2), .I2(n5312), .I3(n5310), 
            .O(n5907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__8454.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__8455 (.I0(n5906), .I1(n5311), .I2(n5313), .I3(n5907), 
            .O(n18593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8455.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8456 (.I0(n4767), .I1(n5330), .O(n5908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8456.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8457 (.I0(\XI[31][16] ), .I1(n5908), .I2(n5334), .I3(n5335), 
            .O(n18592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8457.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8458 (.I0(n4767), .I1(n5336), .I2(MEM_STORE), .I3(STAGE4_EN), 
            .O(ceg_net51753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8458.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8459 (.I0(\XI[31][17] ), .I1(n5908), .I2(n5338), .I3(n5339), 
            .O(n18591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8459.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8460 (.I0(\XI[31][18] ), .I1(n5908), .I2(n5341), .I3(n5342), 
            .O(n18590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8460.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8461 (.I0(\XI[31][19] ), .I1(n5908), .I2(n5344), .I3(n5345), 
            .O(n18589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8461.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8462 (.I0(\XI[31][20] ), .I1(n5908), .I2(n5347), .I3(n5348), 
            .O(n18588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8462.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8463 (.I0(\XI[31][21] ), .I1(n5908), .I2(n5350), .I3(n5351), 
            .O(n18587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8463.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8464 (.I0(\XI[31][22] ), .I1(n5908), .I2(n5353), .I3(n5354), 
            .O(n18586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8464.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8465 (.I0(\XI[31][23] ), .I1(n5908), .I2(n5356), .I3(n5357), 
            .O(n18585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8465.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8466 (.I0(\XI[31][24] ), .I1(n5908), .I2(n5359), .I3(n5360), 
            .O(n18584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8466.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8467 (.I0(\XI[31][25] ), .I1(n5908), .I2(n5362), .I3(n5363), 
            .O(n18583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8467.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8468 (.I0(\XI[31][26] ), .I1(n5908), .I2(n5365), .I3(n5366), 
            .O(n18582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8468.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8469 (.I0(\XI[31][27] ), .I1(n5908), .I2(n5368), .I3(n5369), 
            .O(n18581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8469.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8470 (.I0(\XI[31][28] ), .I1(n5908), .I2(n5371), .I3(n5372), 
            .O(n18580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8470.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8471 (.I0(\XI[31][29] ), .I1(n5908), .I2(n5374), .I3(n5375), 
            .O(n18579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8471.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8472 (.I0(\XI[31][30] ), .I1(n5908), .I2(n5377), .I3(n5378), 
            .O(n18578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8472.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8473 (.I0(\XI[31][31] ), .I1(n5908), .I2(n5380), .I3(n5381), 
            .O(n18577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__8473.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__8474 (.I0(\LOAD_DATA[1] ), .I1(\RES[1] ), .I2(LOAD_OP), 
            .O(n19663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8474.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8475 (.I0(\LOAD_DATA[2] ), .I1(\RES[2] ), .I2(LOAD_OP), 
            .O(n19662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8475.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8476 (.I0(\LOAD_DATA[3] ), .I1(n1612), .I2(LOAD_OP), 
            .O(n19661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8476.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8477 (.I0(\LOAD_DATA[4] ), .I1(n1611), .I2(LOAD_OP), 
            .O(n19660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8477.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8478 (.I0(\LOAD_DATA[5] ), .I1(n1610), .I2(LOAD_OP), 
            .O(n19659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8478.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8479 (.I0(\LOAD_DATA[6] ), .I1(n1609), .I2(LOAD_OP), 
            .O(n19658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8479.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8480 (.I0(\LOAD_DATA[7] ), .I1(n1608), .I2(LOAD_OP), 
            .O(n19657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8480.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8481 (.I0(n2741), .I1(\ARG2[30] ), .I2(\ARG1[30] ), 
            .O(n2738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8481.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8482 (.I0(n3481), .I1(n3472), .I2(n3491), .I3(n3499), 
            .O(n2750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8482.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8483 (.I0(\ARG1[28] ), .I1(\ARG2[28] ), .I2(\ARG2[27] ), 
            .I3(\ARG1[27] ), .O(n5909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__8483.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__8484 (.I0(n2750), .I1(n3500), .I2(n5909), .O(n2744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__8484.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__8485 (.I0(n2750), .I1(\ARG2[27] ), .I2(\ARG1[27] ), 
            .O(n2747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8485.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8486 (.I0(n3481), .I1(n3472), .I2(n3490), .I3(n3496), 
            .O(n5910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8486.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8487 (.I0(n5910), .I1(n3486), .I2(n3487), .I3(n3497), 
            .O(n2753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__8487.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__8488 (.I0(\ARG2[24] ), .I1(\ARG1[24] ), .I2(n5910), 
            .I3(n3486), .O(n2756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__8488.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__8489 (.I0(n5910), .I1(n3486), .O(n2759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__8489.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__8490 (.I0(n3481), .I1(n3472), .I2(n3490), .O(n5911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8490.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8491 (.I0(\ARG2[21] ), .I1(\ARG1[21] ), .I2(n3495), 
            .O(n5912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__8491.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__8492 (.I0(n3482), .I1(n3483), .O(n5913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8492.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8493 (.I0(\ARG1[22] ), .I1(\ARG2[22] ), .O(n5914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8493.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8494 (.I0(n5911), .I1(n5912), .I2(n5913), .I3(n5914), 
            .O(n2762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8494.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8495 (.I0(n5911), .I1(n5912), .I2(n3483), .O(n2765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__8495.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__8496 (.I0(n5911), .I1(n3495), .I2(\ARG2[20] ), .I3(\ARG1[20] ), 
            .O(n2768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__8496.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__8497 (.I0(\ARG2[19] ), .I1(\ARG1[19] ), .I2(n5911), 
            .O(n2771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__8497.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__8498 (.I0(n3481), .I1(n3472), .I2(n3489), .O(n2774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__8498.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__8499 (.I0(n3466), .I1(n3455), .O(n2792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__8499.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__8500 (.I0(n3477), .I1(n3476), .I2(n3480), .O(n5915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__8500.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__8501 (.I0(n2792), .I1(n3471), .I2(n5915), .O(n5916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__8501.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__8502 (.I0(\ARG2[17] ), .I1(n5916), .I2(\ARG1[17] ), 
            .I3(n3467), .O(n2777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7150 */ ;
    defparam LUT__8502.LUTMASK = 16'h7150;
    EFX_LUT4 LUT__8503 (.I0(n5916), .I1(n3467), .O(n2780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8503.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8504 (.I0(\ARG2[13] ), .I1(\ARG1[13] ), .I2(n3466), 
            .I3(n3455), .O(n2789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__8504.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__8505 (.I0(n2789), .I1(\ARG2[14] ), .I2(\ARG1[14] ), 
            .O(n2786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8505.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8506 (.I0(n2786), .I1(\ARG2[15] ), .I2(\ARG1[15] ), 
            .O(n2783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8506.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8507 (.I0(n3477), .I1(n3452), .I2(n3453), .O(n2798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__8507.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__8508 (.I0(n2798), .I1(\ARG2[11] ), .I2(\ARG1[11] ), 
            .O(n2795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8508.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8509 (.I0(n3456), .I1(n3457), .I2(n3459), .O(n5917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8509.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8510 (.I0(n3461), .I1(\ARG2[3] ), .I2(\ARG1[3] ), .I3(n5917), 
            .O(n2819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__8510.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__8511 (.I0(\ARG2[6] ), .I1(\ARG1[6] ), .O(n5918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8511.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8512 (.I0(n2819), .I1(n3458), .I2(n3464), .I3(n5918), 
            .O(n5919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__8512.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__8513 (.I0(\ARG2[7] ), .I1(n3463), .I2(n5919), .I3(\ARG1[7] ), 
            .O(n2807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5701 */ ;
    defparam LUT__8513.LUTMASK = 16'h5701;
    EFX_LUT4 LUT__8514 (.I0(\ARG2[9] ), .I1(\ARG1[9] ), .I2(\ARG1[8] ), 
            .I3(\ARG2[8] ), .O(n5920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__8514.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__8515 (.I0(n2807), .I1(n3451), .I2(n5920), .O(n2801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__8515.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__8516 (.I0(n2807), .I1(\ARG2[8] ), .I2(\ARG1[8] ), .O(n2804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8516.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8517 (.I0(n5919), .I1(n3463), .O(n2810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8517.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8518 (.I0(n2819), .I1(n3458), .I2(n3464), .O(n2813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__8518.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__8519 (.I0(n2819), .I1(\ARG2[4] ), .I2(\ARG1[4] ), .O(n2816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8519.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8520 (.I0(n3456), .I1(n3457), .O(n2825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__8520.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__8521 (.I0(n2825), .I1(\ARG2[2] ), .I2(\ARG1[2] ), .O(n2822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__8521.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__8556 (.I0(\PC[0] ), .O(\PC[0]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__8556.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__8558 (.I0(RST), .O(n1795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__8558.LUTMASK = 16'h5555;
    EFX_LUT4 \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_rtinv  (.I0(\RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_q_pinv ), 
            .O(\RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_rtinv .LUTMASK = 16'h5555;
    EFX_LUT4 \CutToMuxOpt_3/Lut_1  (.I0(\XII[0][5] ), .I1(\XII[1][5] ), 
            .I2(n2953), .I3(\CutToMuxOpt_3/n7 ), .O(n3107)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_3/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_3/Lut_0  (.I0(\XII[2][5] ), .I1(\XII[3][5] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_3/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_3/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_2/Lut_1  (.I0(\XII[8][3] ), .I1(\XII[9][3] ), 
            .I2(n2953), .I3(\CutToMuxOpt_2/n7 ), .O(n3041)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_2/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_2/Lut_0  (.I0(\XII[10][3] ), .I1(\XII[11][3] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_2/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_2/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_1/Lut_1  (.I0(\XII[12][4] ), .I1(\XII[14][4] ), 
            .I2(n2954), .I3(\CutToMuxOpt_1/n7 ), .O(n3013)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_1/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_1/Lut_0  (.I0(\XII[13][4] ), .I1(\XII[15][4] ), 
            .I2(n2954), .I3(n51766), .O(\CutToMuxOpt_1/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_1/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_0/Lut_1  (.I0(\XII[8][4] ), .I1(\XII[10][4] ), 
            .I2(n2954), .I3(\CutToMuxOpt_0/n7 ), .O(n3010)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_0/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_0/Lut_0  (.I0(\XII[9][4] ), .I1(\XII[11][4] ), 
            .I2(n2954), .I3(n51766), .O(\CutToMuxOpt_0/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_0/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_23/Lut_1  (.I0(\XI[0][22] ), .I1(\XI[1][22] ), 
            .I2(n2953), .I3(\CutToMuxOpt_23/n7 ), .O(n3937)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_23/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_23/Lut_0  (.I0(\XI[2][22] ), .I1(\XI[3][22] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_23/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_23/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_22/Lut_1  (.I0(\XI[0][30] ), .I1(\XI[1][30] ), 
            .I2(n2953), .I3(\CutToMuxOpt_22/n7 ), .O(n3882)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_22/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_22/Lut_0  (.I0(\XI[2][30] ), .I1(\XI[3][30] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_22/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_22/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_21/Lut_1  (.I0(\XI[0][23] ), .I1(\XI[1][23] ), 
            .I2(n2953), .I3(\CutToMuxOpt_21/n7 ), .O(n3852)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_21/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_21/Lut_0  (.I0(\XI[2][23] ), .I1(\XI[3][23] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_21/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_21/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_20/Lut_1  (.I0(\XI[0][31] ), .I1(\XI[1][31] ), 
            .I2(n2953), .I3(\CutToMuxOpt_20/n7 ), .O(n3822)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_20/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_20/Lut_0  (.I0(\XI[2][31] ), .I1(\XI[3][31] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_20/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_20/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_19/Lut_1  (.I0(\XI[0][24] ), .I1(\XI[1][24] ), 
            .I2(n2953), .I3(\CutToMuxOpt_19/n7 ), .O(n3792)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_19/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_19/Lut_0  (.I0(\XI[2][24] ), .I1(\XI[3][24] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_19/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_19/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_18/Lut_1  (.I0(\XI[0][25] ), .I1(\XI[1][25] ), 
            .I2(n2953), .I3(\CutToMuxOpt_18/n7 ), .O(n3762)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_18/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_18/Lut_0  (.I0(\XI[2][25] ), .I1(\XI[3][25] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_18/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_18/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_17/Lut_1  (.I0(\XI[0][19] ), .I1(\XI[1][19] ), 
            .I2(n2953), .I3(\CutToMuxOpt_17/n7 ), .O(n3732)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_17/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_17/Lut_0  (.I0(\XI[2][19] ), .I1(\XI[3][19] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_17/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_17/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_16/Lut_1  (.I0(\XI[0][18] ), .I1(\XI[1][18] ), 
            .I2(n2953), .I3(\CutToMuxOpt_16/n7 ), .O(n3702)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_16/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_16/Lut_0  (.I0(\XI[2][18] ), .I1(\XI[3][18] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_16/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_16/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_15/Lut_1  (.I0(\XI[0][17] ), .I1(\XI[1][17] ), 
            .I2(n2953), .I3(\CutToMuxOpt_15/n7 ), .O(n3672)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_15/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_15/Lut_0  (.I0(\XI[2][17] ), .I1(\XI[3][17] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_15/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_15/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_14/Lut_1  (.I0(\XI[0][16] ), .I1(\XI[1][16] ), 
            .I2(n2953), .I3(\CutToMuxOpt_14/n7 ), .O(n3642)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_14/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_14/Lut_0  (.I0(\XI[2][16] ), .I1(\XI[3][16] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_14/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_14/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_13/Lut_1  (.I0(\XI[0][15] ), .I1(\XI[1][15] ), 
            .I2(n2953), .I3(\CutToMuxOpt_13/n7 ), .O(n3612)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_13/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_13/Lut_0  (.I0(\XI[2][15] ), .I1(\XI[3][15] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_13/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_13/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \CutToMuxOpt_12/Lut_1  (.I0(\XI[0][14] ), .I1(\XI[1][14] ), 
            .I2(n2953), .I3(\CutToMuxOpt_12/n7 ), .O(n3582)) /* verific LUTMASK=16'hf305, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_12/Lut_1 .LUTMASK = 16'hf305;
    EFX_LUT4 \CutToMuxOpt_12/Lut_0  (.I0(\XI[2][14] ), .I1(\XI[3][14] ), 
            .I2(n2953), .I3(n51770), .O(\CutToMuxOpt_12/n7 )) /* verific LUTMASK=16'h3f50, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4 */ ;
    defparam \CutToMuxOpt_12/Lut_0 .LUTMASK = 16'h3f50;
    EFX_LUT4 \RES[22]_2~FF_brt_41_brt_97_brt_168_rtinv  (.I0(\RES[22]_2~FF_brt_41_brt_97_brt_168_q_pinv ), 
            .O(\RES[22]_2~FF_brt_41_brt_97_brt_168_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168_rtinv .LUTMASK = 16'h5555;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(CLK), .O(\CLK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i3  (.I0(n2825), .I1(1'b1), .CI(1'b0), 
            .CO(n5951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i4  (.I0(n2822), .I1(1'b1), .CI(1'b0), 
            .CO(n5950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i5  (.I0(n2819), .I1(1'b1), .CI(1'b0), 
            .CO(n5949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i6  (.I0(n2816), .I1(1'b1), .CI(1'b0), 
            .CO(n5948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i7  (.I0(n2813), .I1(1'b1), .CI(1'b0), 
            .CO(n5947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i8  (.I0(n2810), .I1(1'b1), .CI(1'b0), 
            .CO(n5946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i9  (.I0(n2807), .I1(1'b1), .CI(1'b0), 
            .CO(n5945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i10  (.I0(n2804), .I1(1'b1), .CI(1'b0), 
            .CO(n5944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i11  (.I0(n2801), .I1(1'b1), .CI(1'b0), 
            .CO(n5943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i12  (.I0(n2798), .I1(1'b1), .CI(1'b0), 
            .CO(n5942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i13  (.I0(n2795), .I1(1'b1), .CI(1'b0), 
            .CO(n5941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i14  (.I0(n2792), .I1(1'b1), .CI(1'b0), 
            .CO(n5940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i15  (.I0(n2789), .I1(1'b1), .CI(1'b0), 
            .CO(n5939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i16  (.I0(n2786), .I1(1'b1), .CI(1'b0), 
            .CO(n5938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i17  (.I0(n2783), .I1(1'b1), .CI(1'b0), 
            .CO(n5937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i18  (.I0(n2780), .I1(1'b1), .CI(1'b0), 
            .CO(n5936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i19  (.I0(n2777), .I1(1'b1), .CI(1'b0), 
            .CO(n5935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i20  (.I0(n2774), .I1(1'b1), .CI(1'b0), 
            .CO(n5934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i21  (.I0(n2771), .I1(1'b1), .CI(1'b0), 
            .CO(n5933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i22  (.I0(n2768), .I1(1'b1), .CI(1'b0), 
            .CO(n5932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i23  (.I0(n2765), .I1(1'b1), .CI(1'b0), 
            .CO(n5931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i24  (.I0(n2762), .I1(1'b1), .CI(1'b0), 
            .CO(n5930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i25  (.I0(n2759), .I1(1'b1), .CI(1'b0), 
            .CO(n5929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i25 .I1_POLARITY = 1'b1;
    EFX_FF \RES[31]_2~FF_brt_66_brt_119_brt_191  (.D(n1341), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[31]_2~FF_brt_66_brt_119_brt_191_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191 .CLK_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191 .CE_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191 .SR_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191 .D_POLARITY = 1'b0;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191 .SR_SYNC = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191 .SR_VALUE = 1'b0;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[31]_2~FF_brt_66_brt_119_brt_190  (.D(n1389), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[31]_2~FF_brt_66_brt_119_brt_190_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_190 .CLK_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_190 .CE_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_190 .SR_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_190 .D_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_190 .SR_SYNC = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_190 .SR_VALUE = 1'b0;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_190 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[30]_2~FF_brt_189  (.D(n5299), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[30]_2~FF_brt_189_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[30]_2~FF_brt_189 .CLK_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_189 .CE_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_189 .SR_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_189 .D_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_189 .SR_SYNC = 1'b1;
    defparam \RES[30]_2~FF_brt_189 .SR_VALUE = 1'b0;
    defparam \RES[30]_2~FF_brt_189 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[30]_2~FF_brt_188  (.D(n5297), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[30]_2~FF_brt_188_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[30]_2~FF_brt_188 .CLK_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_188 .CE_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_188 .SR_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_188 .D_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_188 .SR_SYNC = 1'b1;
    defparam \RES[30]_2~FF_brt_188 .SR_VALUE = 1'b0;
    defparam \RES[30]_2~FF_brt_188 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[30]_2~FF_brt_187  (.D(n5294), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[30]_2~FF_brt_187_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[30]_2~FF_brt_187 .CLK_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_187 .CE_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_187 .SR_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_187 .D_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_187 .SR_SYNC = 1'b1;
    defparam \RES[30]_2~FF_brt_187 .SR_VALUE = 1'b0;
    defparam \RES[30]_2~FF_brt_187 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[30]_2~FF_brt_186  (.D(n5295), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[30]_2~FF_brt_186_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[30]_2~FF_brt_186 .CLK_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_186 .CE_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_186 .SR_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_186 .D_POLARITY = 1'b1;
    defparam \RES[30]_2~FF_brt_186 .SR_SYNC = 1'b1;
    defparam \RES[30]_2~FF_brt_186 .SR_VALUE = 1'b0;
    defparam \RES[30]_2~FF_brt_186 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185  (.D(n1392), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185 .CLK_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185 .CE_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185 .SR_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185 .D_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185 .SR_SYNC = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185 .SR_VALUE = 1'b0;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_185 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184  (.D(n1343), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184 .CLK_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184 .CE_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184 .SR_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184 .D_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184 .SR_SYNC = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184 .SR_VALUE = 1'b0;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_117_brt_184 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183  (.D(n1394), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183 .D_POLARITY = 1'b0;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_183 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182  (.D(n1344), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182 .D_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_115_brt_182 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[27]_2~FF_brt_55_brt_113_brt_181  (.D(n5264), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[27]_2~FF_brt_55_brt_113_brt_181_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_181 .CLK_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_181 .CE_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_181 .SR_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_181 .D_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_181 .SR_SYNC = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_181 .SR_VALUE = 1'b0;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_181 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[27]_2~FF_brt_55_brt_113_brt_180  (.D(n5263), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[27]_2~FF_brt_55_brt_113_brt_180_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_180 .CLK_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_180 .CE_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_180 .SR_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_180 .D_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_180 .SR_SYNC = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_180 .SR_VALUE = 1'b0;
    defparam \RES[27]_2~FF_brt_55_brt_113_brt_180 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179  (.D(n1398), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179 .CLK_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179 .CE_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179 .SR_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179 .D_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179 .SR_SYNC = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179 .SR_VALUE = 1'b0;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_179 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178  (.D(n1346), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178 .CLK_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178 .CE_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178 .SR_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178 .D_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178 .SR_SYNC = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178 .SR_VALUE = 1'b0;
    defparam \RES[26]_2~FF_brt_10_brt_52_brt_110_brt_178 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[25]_2~FF_brt_108_brt_177  (.D(n5243), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[25]_2~FF_brt_108_brt_177_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[25]_2~FF_brt_108_brt_177 .CLK_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_177 .CE_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_177 .SR_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_177 .D_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_177 .SR_SYNC = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_177 .SR_VALUE = 1'b0;
    defparam \RES[25]_2~FF_brt_108_brt_177 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[25]_2~FF_brt_108_brt_176  (.D(n5242), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[25]_2~FF_brt_108_brt_176_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[25]_2~FF_brt_108_brt_176 .CLK_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_176 .CE_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_176 .SR_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_176 .D_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_176 .SR_SYNC = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_176 .SR_VALUE = 1'b0;
    defparam \RES[25]_2~FF_brt_108_brt_176 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[25]_2~FF_brt_108_brt_175  (.D(n1347), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[25]_2~FF_brt_108_brt_175_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[25]_2~FF_brt_108_brt_175 .CLK_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_175 .CE_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_175 .SR_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_175 .D_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_175 .SR_SYNC = 1'b1;
    defparam \RES[25]_2~FF_brt_108_brt_175 .SR_VALUE = 1'b0;
    defparam \RES[25]_2~FF_brt_108_brt_175 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_49_brt_105_brt_174  (.D(n5233), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[24]_2~FF_brt_49_brt_105_brt_174_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_174 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_174 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_174 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_174 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_174 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_174 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_174 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_49_brt_105_brt_173  (.D(n1348), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[24]_2~FF_brt_49_brt_105_brt_173_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_173 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_173 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_173 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_173 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_173 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_173 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_173 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_49_brt_105_brt_172  (.D(n5232), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[24]_2~FF_brt_49_brt_105_brt_172_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_172 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_172 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_172 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_172 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_172 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_172 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_49_brt_105_brt_172 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[23]_2~FF_brt_45_brt_99_brt_171  (.D(n1349), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[23]_2~FF_brt_45_brt_99_brt_171_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_171 .CLK_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_171 .CE_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_171 .SR_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_171 .D_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_171 .SR_SYNC = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_171 .SR_VALUE = 1'b0;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_171 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[23]_2~FF_brt_45_brt_99_brt_170  (.D(n1404), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[23]_2~FF_brt_45_brt_99_brt_170_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_170 .CLK_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_170 .CE_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_170 .SR_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_170 .D_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_170 .SR_SYNC = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_170 .SR_VALUE = 1'b0;
    defparam \RES[23]_2~FF_brt_45_brt_99_brt_170 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[22]_2~FF_brt_41_brt_97_brt_169  (.D(n5166), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[22]_2~FF_brt_41_brt_97_brt_169_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_169 .CLK_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_169 .CE_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_169 .SR_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_169 .D_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_169 .SR_SYNC = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_169 .SR_VALUE = 1'b0;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_169 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[22]_2~FF_brt_41_brt_97_brt_168  (.D(n1350), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[22]_2~FF_brt_41_brt_97_brt_168_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168 .CLK_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168 .CE_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168 .SR_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168 .D_POLARITY = 1'b0;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168 .SR_SYNC = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168 .SR_VALUE = 1'b0;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_168 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[22]_2~FF_brt_41_brt_97_brt_167  (.D(n1406), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[22]_2~FF_brt_41_brt_97_brt_167_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_167 .CLK_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_167 .CE_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_167 .SR_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_167 .D_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_167 .SR_SYNC = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_167 .SR_VALUE = 1'b0;
    defparam \RES[22]_2~FF_brt_41_brt_97_brt_167 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[21]_2~FF_brt_96_brt_166  (.D(n1408), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[21]_2~FF_brt_96_brt_166_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[21]_2~FF_brt_96_brt_166 .CLK_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_166 .CE_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_166 .SR_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_166 .D_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_166 .SR_SYNC = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_166 .SR_VALUE = 1'b0;
    defparam \RES[21]_2~FF_brt_96_brt_166 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[21]_2~FF_brt_96_brt_165  (.D(n1351), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[21]_2~FF_brt_96_brt_165_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[21]_2~FF_brt_96_brt_165 .CLK_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_165 .CE_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_165 .SR_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_165 .D_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_165 .SR_SYNC = 1'b1;
    defparam \RES[21]_2~FF_brt_96_brt_165 .SR_VALUE = 1'b0;
    defparam \RES[21]_2~FF_brt_96_brt_165 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[20]_2~FF_brt_93_brt_164  (.D(n3552), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[20]_2~FF_brt_93_brt_164_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[20]_2~FF_brt_93_brt_164 .CLK_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_164 .CE_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_164 .SR_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_164 .D_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_164 .SR_SYNC = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_164 .SR_VALUE = 1'b0;
    defparam \RES[20]_2~FF_brt_93_brt_164 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[20]_2~FF_brt_93_brt_163  (.D(n1410), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[20]_2~FF_brt_93_brt_163_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[20]_2~FF_brt_93_brt_163 .CLK_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_163 .CE_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_163 .SR_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_163 .D_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_163 .SR_SYNC = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_163 .SR_VALUE = 1'b0;
    defparam \RES[20]_2~FF_brt_93_brt_163 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[20]_2~FF_brt_93_brt_162  (.D(n1352), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[20]_2~FF_brt_93_brt_162_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[20]_2~FF_brt_93_brt_162 .CLK_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_162 .CE_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_162 .SR_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_162 .D_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_162 .SR_SYNC = 1'b1;
    defparam \RES[20]_2~FF_brt_93_brt_162 .SR_VALUE = 1'b0;
    defparam \RES[20]_2~FF_brt_93_brt_162 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[19]_2~FF_brt_161  (.D(n5181), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[19]_2~FF_brt_161_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[19]_2~FF_brt_161 .CLK_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_161 .CE_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_161 .SR_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_161 .D_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_161 .SR_SYNC = 1'b1;
    defparam \RES[19]_2~FF_brt_161 .SR_VALUE = 1'b0;
    defparam \RES[19]_2~FF_brt_161 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[19]_2~FF_brt_160  (.D(n5180), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[19]_2~FF_brt_160_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[19]_2~FF_brt_160 .CLK_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_160 .CE_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_160 .SR_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_160 .D_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_160 .SR_SYNC = 1'b1;
    defparam \RES[19]_2~FF_brt_160 .SR_VALUE = 1'b0;
    defparam \RES[19]_2~FF_brt_160 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[19]_2~FF_brt_159  (.D(n5178), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[19]_2~FF_brt_159_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[19]_2~FF_brt_159 .CLK_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_159 .CE_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_159 .SR_POLARITY = 1'b1;
    defparam \RES[19]_2~FF_brt_159 .D_POLARITY = 1'b0;
    defparam \RES[19]_2~FF_brt_159 .SR_SYNC = 1'b1;
    defparam \RES[19]_2~FF_brt_159 .SR_VALUE = 1'b0;
    defparam \RES[19]_2~FF_brt_159 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[18]_2~FF_brt_90_brt_157  (.D(n1414), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[18]_2~FF_brt_90_brt_157_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[18]_2~FF_brt_90_brt_157 .CLK_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_157 .CE_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_157 .SR_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_157 .D_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_157 .SR_SYNC = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_157 .SR_VALUE = 1'b0;
    defparam \RES[18]_2~FF_brt_90_brt_157 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[18]_2~FF_brt_90_brt_156  (.D(n1354), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[18]_2~FF_brt_90_brt_156_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[18]_2~FF_brt_90_brt_156 .CLK_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_156 .CE_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_156 .SR_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_156 .D_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_156 .SR_SYNC = 1'b1;
    defparam \RES[18]_2~FF_brt_90_brt_156 .SR_VALUE = 1'b0;
    defparam \RES[18]_2~FF_brt_90_brt_156 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155  (.D(n1416), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_155 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154  (.D(n1355), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_87_brt_154 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153  (.D(n1418), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153 .CLK_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153 .CE_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153 .SR_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153 .D_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153 .SR_SYNC = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153 .SR_VALUE = 1'b0;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_153 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152  (.D(n1356), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152 .CLK_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152 .CE_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152 .SR_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152 .D_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152 .SR_SYNC = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152 .SR_VALUE = 1'b0;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_84_brt_152 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[15]_2~FF_brt_30_brt_82_brt_151  (.D(n5128), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[15]_2~FF_brt_30_brt_82_brt_151_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151 .CLK_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151 .CE_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151 .SR_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151 .D_POLARITY = 1'b0;
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151 .SR_SYNC = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151 .SR_VALUE = 1'b0;
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[14]_2~FF_brt_150  (.D(n5119), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[14]_2~FF_brt_150_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[14]_2~FF_brt_150 .CLK_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_150 .CE_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_150 .SR_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_150 .D_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_150 .SR_SYNC = 1'b1;
    defparam \RES[14]_2~FF_brt_150 .SR_VALUE = 1'b0;
    defparam \RES[14]_2~FF_brt_150 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[14]_2~FF_brt_149  (.D(n5116), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[14]_2~FF_brt_149_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[14]_2~FF_brt_149 .CLK_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_149 .CE_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_149 .SR_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_149 .D_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_149 .SR_SYNC = 1'b1;
    defparam \RES[14]_2~FF_brt_149 .SR_VALUE = 1'b0;
    defparam \RES[14]_2~FF_brt_149 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[14]_2~FF_brt_148  (.D(n5110), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[14]_2~FF_brt_148_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[14]_2~FF_brt_148 .CLK_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_148 .CE_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_148 .SR_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_148 .D_POLARITY = 1'b1;
    defparam \RES[14]_2~FF_brt_148 .SR_SYNC = 1'b1;
    defparam \RES[14]_2~FF_brt_148 .SR_VALUE = 1'b0;
    defparam \RES[14]_2~FF_brt_148 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[13]_2~FF_brt_147  (.D(n5099), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[13]_2~FF_brt_147_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[13]_2~FF_brt_147 .CLK_POLARITY = 1'b1;
    defparam \RES[13]_2~FF_brt_147 .CE_POLARITY = 1'b1;
    defparam \RES[13]_2~FF_brt_147 .SR_POLARITY = 1'b1;
    defparam \RES[13]_2~FF_brt_147 .D_POLARITY = 1'b0;
    defparam \RES[13]_2~FF_brt_147 .SR_SYNC = 1'b1;
    defparam \RES[13]_2~FF_brt_147 .SR_VALUE = 1'b0;
    defparam \RES[13]_2~FF_brt_147 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[13]_2~FF_brt_146  (.D(n5105), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[13]_2~FF_brt_146_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[13]_2~FF_brt_146 .CLK_POLARITY = 1'b1;
    defparam \RES[13]_2~FF_brt_146 .CE_POLARITY = 1'b1;
    defparam \RES[13]_2~FF_brt_146 .SR_POLARITY = 1'b1;
    defparam \RES[13]_2~FF_brt_146 .D_POLARITY = 1'b0;
    defparam \RES[13]_2~FF_brt_146 .SR_SYNC = 1'b1;
    defparam \RES[13]_2~FF_brt_146 .SR_VALUE = 1'b0;
    defparam \RES[13]_2~FF_brt_146 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[12]_2~FF_brt_78_brt_145  (.D(n5084), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[12]_2~FF_brt_78_brt_145_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[12]_2~FF_brt_78_brt_145 .CLK_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_78_brt_145 .CE_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_78_brt_145 .SR_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_78_brt_145 .D_POLARITY = 1'b0;
    defparam \RES[12]_2~FF_brt_78_brt_145 .SR_SYNC = 1'b1;
    defparam \RES[12]_2~FF_brt_78_brt_145 .SR_VALUE = 1'b0;
    defparam \RES[12]_2~FF_brt_78_brt_145 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[11]_2~FF_brt_144  (.D(n5079), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[11]_2~FF_brt_144_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[11]_2~FF_brt_144 .CLK_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_144 .CE_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_144 .SR_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_144 .D_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_144 .SR_SYNC = 1'b1;
    defparam \RES[11]_2~FF_brt_144 .SR_VALUE = 1'b0;
    defparam \RES[11]_2~FF_brt_144 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[11]_2~FF_brt_143  (.D(n5077), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[11]_2~FF_brt_143_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[11]_2~FF_brt_143 .CLK_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_143 .CE_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_143 .SR_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_143 .D_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_143 .SR_SYNC = 1'b1;
    defparam \RES[11]_2~FF_brt_143 .SR_VALUE = 1'b0;
    defparam \RES[11]_2~FF_brt_143 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[11]_2~FF_brt_142  (.D(n5068), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[11]_2~FF_brt_142_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[11]_2~FF_brt_142 .CLK_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_142 .CE_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_142 .SR_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_142 .D_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_142 .SR_SYNC = 1'b1;
    defparam \RES[11]_2~FF_brt_142 .SR_VALUE = 1'b0;
    defparam \RES[11]_2~FF_brt_142 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[11]_2~FF_brt_141  (.D(n5074), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[11]_2~FF_brt_141_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[11]_2~FF_brt_141 .CLK_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_141 .CE_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_141 .SR_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_141 .D_POLARITY = 1'b1;
    defparam \RES[11]_2~FF_brt_141 .SR_SYNC = 1'b1;
    defparam \RES[11]_2~FF_brt_141 .SR_VALUE = 1'b0;
    defparam \RES[11]_2~FF_brt_141 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140  (.D(n1430), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140 .CLK_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140 .CE_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140 .SR_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140 .D_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140 .SR_SYNC = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140 .SR_VALUE = 1'b0;
    defparam \RES[10]_2~FF_brt_3_brt_28_brt_76_brt_140 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[0]_2~FF_brt_192  (.D(n3540), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[0]_2~FF_brt_192_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[0]_2~FF_brt_192 .CLK_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_192 .CE_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_192 .SR_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_192 .D_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_192 .SR_SYNC = 1'b1;
    defparam \RES[0]_2~FF_brt_192 .SR_VALUE = 1'b0;
    defparam \RES[0]_2~FF_brt_192 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[31]_2~FF_brt_66_brt_118  (.D(\ARG1[31] ), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[31]_2~FF_brt_66_brt_118_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[31]_2~FF_brt_66_brt_118 .CLK_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_118 .CE_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_118 .SR_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_118 .D_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_118 .SR_SYNC = 1'b1;
    defparam \RES[31]_2~FF_brt_66_brt_118 .SR_VALUE = 1'b0;
    defparam \RES[31]_2~FF_brt_66_brt_118 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[0]_2~FF_brt_194  (.D(n2741), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[0]_2~FF_brt_194_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[0]_2~FF_brt_194 .CLK_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_194 .CE_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_194 .SR_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_194 .D_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_194 .SR_SYNC = 1'b1;
    defparam \RES[0]_2~FF_brt_194 .SR_VALUE = 1'b0;
    defparam \RES[0]_2~FF_brt_194 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[29]_2~FF_brt_16_brt_63_brt_116  (.D(n5284), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[29]_2~FF_brt_16_brt_63_brt_116_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_116 .CLK_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_116 .CE_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_116 .SR_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_116 .D_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_116 .SR_SYNC = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_116 .SR_VALUE = 1'b0;
    defparam \RES[29]_2~FF_brt_16_brt_63_brt_116 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[0]_2~FF_brt_195  (.D(n3504), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[0]_2~FF_brt_195_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[0]_2~FF_brt_195 .CLK_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_195 .CE_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_195 .SR_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_195 .D_POLARITY = 1'b1;
    defparam \RES[0]_2~FF_brt_195 .SR_SYNC = 1'b1;
    defparam \RES[0]_2~FF_brt_195 .SR_VALUE = 1'b0;
    defparam \RES[0]_2~FF_brt_195 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_15_brt_60_brt_114  (.D(n5269), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[28]_2~FF_brt_15_brt_60_brt_114_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_114 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_114 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_114 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_114 .D_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_114 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_114 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_15_brt_60_brt_114 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[19]_2~FF_brt_159_rtinv  (.I0(\RES[19]_2~FF_brt_159_q_pinv ), 
            .O(\RES[19]_2~FF_brt_159_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[19]_2~FF_brt_159_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[27]_2~FF_brt_55_brt_112  (.D(n5259), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[27]_2~FF_brt_55_brt_112_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[27]_2~FF_brt_55_brt_112 .CLK_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_112 .CE_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_112 .SR_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_112 .D_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_112 .SR_SYNC = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_112 .SR_VALUE = 1'b0;
    defparam \RES[27]_2~FF_brt_55_brt_112 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[27]_2~FF_brt_55_brt_111  (.D(n5262), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[27]_2~FF_brt_55_brt_111_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[27]_2~FF_brt_55_brt_111 .CLK_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_111 .CE_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_111 .SR_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_111 .D_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_111 .SR_SYNC = 1'b1;
    defparam \RES[27]_2~FF_brt_55_brt_111 .SR_VALUE = 1'b0;
    defparam \RES[27]_2~FF_brt_55_brt_111 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[15]_2~FF_brt_30_brt_82_brt_151_rtinv  (.I0(\RES[15]_2~FF_brt_30_brt_82_brt_151_q_pinv ), 
            .O(\RES[15]_2~FF_brt_30_brt_82_brt_151_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[15]_2~FF_brt_30_brt_82_brt_151_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[25]_2~FF_brt_109  (.D(n5247), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[25]_2~FF_brt_109_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[25]_2~FF_brt_109 .CLK_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_109 .CE_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_109 .SR_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_109 .D_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_109 .SR_SYNC = 1'b1;
    defparam \RES[25]_2~FF_brt_109 .SR_VALUE = 1'b0;
    defparam \RES[25]_2~FF_brt_109 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[13]_2~FF_brt_147_rtinv  (.I0(\RES[13]_2~FF_brt_147_q_pinv ), 
            .O(\RES[13]_2~FF_brt_147_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[13]_2~FF_brt_147_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[25]_2~FF_brt_107  (.D(n5240), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[25]_2~FF_brt_107_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[25]_2~FF_brt_107 .CLK_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_107 .CE_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_107 .SR_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_107 .D_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_107 .SR_SYNC = 1'b1;
    defparam \RES[25]_2~FF_brt_107 .SR_VALUE = 1'b0;
    defparam \RES[25]_2~FF_brt_107 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[25]_2~FF_brt_106  (.D(n5241), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[25]_2~FF_brt_106_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[25]_2~FF_brt_106 .CLK_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_106 .CE_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_106 .SR_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_106 .D_POLARITY = 1'b1;
    defparam \RES[25]_2~FF_brt_106 .SR_SYNC = 1'b1;
    defparam \RES[25]_2~FF_brt_106 .SR_VALUE = 1'b0;
    defparam \RES[25]_2~FF_brt_106 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[13]_2~FF_brt_146_rtinv  (.I0(\RES[13]_2~FF_brt_146_q_pinv ), 
            .O(\RES[13]_2~FF_brt_146_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[13]_2~FF_brt_146_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[24]_2~FF_brt_49_brt_104  (.D(n5231), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[24]_2~FF_brt_49_brt_104_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_49_brt_104 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_104 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_104 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_104 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_104 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_104 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_49_brt_104 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_49_brt_103  (.D(n5230), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[24]_2~FF_brt_49_brt_103_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_49_brt_103 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_103 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_103 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_103 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_103 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_103 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_49_brt_103 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_49_brt_102  (.D(n5229), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[24]_2~FF_brt_49_brt_102_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_49_brt_102 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_102 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_102 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_102 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_102 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_49_brt_102 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_49_brt_102 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[23]_2~FF_brt_45_brt_100  (.D(n3552), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[23]_2~FF_brt_45_brt_100_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[23]_2~FF_brt_45_brt_100 .CLK_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_100 .CE_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_100 .SR_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_100 .D_POLARITY = 1'b0;
    defparam \RES[23]_2~FF_brt_45_brt_100 .SR_SYNC = 1'b1;
    defparam \RES[23]_2~FF_brt_45_brt_100 .SR_VALUE = 1'b0;
    defparam \RES[23]_2~FF_brt_45_brt_100 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[12]_2~FF_brt_78_brt_145_rtinv  (.I0(\RES[12]_2~FF_brt_78_brt_145_q_pinv ), 
            .O(\RES[12]_2~FF_brt_78_brt_145_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[12]_2~FF_brt_78_brt_145_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[22]_2~FF_brt_41_brt_98  (.D(\OPERATION[3] ), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[22]_2~FF_brt_41_brt_98_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[22]_2~FF_brt_41_brt_98 .CLK_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_98 .CE_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_98 .SR_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_98 .D_POLARITY = 1'b0;
    defparam \RES[22]_2~FF_brt_41_brt_98 .SR_SYNC = 1'b1;
    defparam \RES[22]_2~FF_brt_41_brt_98 .SR_VALUE = 1'b0;
    defparam \RES[22]_2~FF_brt_41_brt_98 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[23]_2~FF_brt_45_brt_100_rtinv  (.I0(\RES[23]_2~FF_brt_45_brt_100_q_pinv ), 
            .O(\RES[23]_2~FF_brt_45_brt_100_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[23]_2~FF_brt_45_brt_100_rtinv .LUTMASK = 16'h5555;
    EFX_LUT4 \RES[20]_2~FF_brt_92_rtinv  (.I0(\RES[20]_2~FF_brt_92_q_pinv ), 
            .O(\RES[20]_2~FF_brt_92_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[20]_2~FF_brt_92_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[21]_2~FF_brt_95  (.D(n5192), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[21]_2~FF_brt_95_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[21]_2~FF_brt_95 .CLK_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_95 .CE_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_95 .SR_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_95 .D_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_95 .SR_SYNC = 1'b1;
    defparam \RES[21]_2~FF_brt_95 .SR_VALUE = 1'b0;
    defparam \RES[21]_2~FF_brt_95 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[21]_2~FF_brt_94  (.D(n5200), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[21]_2~FF_brt_94_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[21]_2~FF_brt_94 .CLK_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_94 .CE_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_94 .SR_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_94 .D_POLARITY = 1'b1;
    defparam \RES[21]_2~FF_brt_94 .SR_SYNC = 1'b1;
    defparam \RES[21]_2~FF_brt_94 .SR_VALUE = 1'b0;
    defparam \RES[21]_2~FF_brt_94 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[18]_2~FF_brt_89_rtinv  (.I0(\RES[18]_2~FF_brt_89_q_pinv ), 
            .O(\RES[18]_2~FF_brt_89_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[18]_2~FF_brt_89_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[20]_2~FF_brt_92  (.D(n5185), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[20]_2~FF_brt_92_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[20]_2~FF_brt_92 .CLK_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_92 .CE_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_92 .SR_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_92 .D_POLARITY = 1'b0;
    defparam \RES[20]_2~FF_brt_92 .SR_SYNC = 1'b1;
    defparam \RES[20]_2~FF_brt_92 .SR_VALUE = 1'b0;
    defparam \RES[20]_2~FF_brt_92 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[20]_2~FF_brt_91  (.D(n5190), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[20]_2~FF_brt_91_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[20]_2~FF_brt_91 .CLK_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_91 .CE_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_91 .SR_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_91 .D_POLARITY = 1'b1;
    defparam \RES[20]_2~FF_brt_91 .SR_SYNC = 1'b1;
    defparam \RES[20]_2~FF_brt_91 .SR_VALUE = 1'b0;
    defparam \RES[20]_2~FF_brt_91 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[3]_2~FF_brt_120_rtinv  (.I0(\RES[3]_2~FF_brt_120_q_pinv ), 
            .O(\RES[3]_2~FF_brt_120_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[3]_2~FF_brt_120_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[18]_2~FF_brt_89  (.D(n5158), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[18]_2~FF_brt_89_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[18]_2~FF_brt_89 .CLK_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_89 .CE_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_89 .SR_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_89 .D_POLARITY = 1'b0;
    defparam \RES[18]_2~FF_brt_89 .SR_SYNC = 1'b1;
    defparam \RES[18]_2~FF_brt_89 .SR_VALUE = 1'b0;
    defparam \RES[18]_2~FF_brt_89 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[18]_2~FF_brt_88  (.D(n5168), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[18]_2~FF_brt_88_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[18]_2~FF_brt_88 .CLK_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_88 .CE_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_88 .SR_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_88 .D_POLARITY = 1'b1;
    defparam \RES[18]_2~FF_brt_88 .SR_SYNC = 1'b1;
    defparam \RES[18]_2~FF_brt_88 .SR_VALUE = 1'b0;
    defparam \RES[18]_2~FF_brt_88 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \RES[31]_2~FF_brt_66_brt_119_brt_191_rtinv  (.I0(\RES[31]_2~FF_brt_66_brt_119_brt_191_q_pinv ), 
            .O(\RES[31]_2~FF_brt_66_brt_119_brt_191_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \RES[31]_2~FF_brt_66_brt_119_brt_191_rtinv .LUTMASK = 16'h5555;
    EFX_FF \RES[17]_2~FF_brt_8_brt_37_brt_86  (.D(n3542), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[17]_2~FF_brt_8_brt_37_brt_86_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_86 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_86 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_86 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_86 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_86 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_86 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_86 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_8_brt_37_brt_85  (.D(n4897), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[17]_2~FF_brt_8_brt_37_brt_85_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_85 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_85 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_85 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_85 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_85 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_85 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_8_brt_37_brt_85 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[16]_2~FF_brt_5_brt_33_brt_83  (.D(n5136), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[16]_2~FF_brt_5_brt_33_brt_83_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_83 .CLK_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_83 .CE_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_83 .SR_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_83 .D_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_83 .SR_SYNC = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_83 .SR_VALUE = 1'b0;
    defparam \RES[16]_2~FF_brt_5_brt_33_brt_83 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[31]_2~FF_brt_67  (.D(n5308), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[31]_2~FF_brt_67_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[31]_2~FF_brt_67 .CLK_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_67 .CE_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_67 .SR_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_67 .D_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_67 .SR_SYNC = 1'b1;
    defparam \RES[31]_2~FF_brt_67 .SR_VALUE = 1'b0;
    defparam \RES[31]_2~FF_brt_67 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[3]_2~FF_brt_120  (.D(n4944), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[3]_2~FF_brt_120_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[3]_2~FF_brt_120 .CLK_POLARITY = 1'b1;
    defparam \RES[3]_2~FF_brt_120 .CE_POLARITY = 1'b1;
    defparam \RES[3]_2~FF_brt_120 .SR_POLARITY = 1'b1;
    defparam \RES[3]_2~FF_brt_120 .D_POLARITY = 1'b0;
    defparam \RES[3]_2~FF_brt_120 .SR_SYNC = 1'b1;
    defparam \RES[3]_2~FF_brt_120 .SR_VALUE = 1'b0;
    defparam \RES[3]_2~FF_brt_120 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[31]_2~FF_brt_65  (.D(n5300), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[31]_2~FF_brt_65_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[31]_2~FF_brt_65 .CLK_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_65 .CE_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_65 .SR_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_65 .D_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_65 .SR_SYNC = 1'b1;
    defparam \RES[31]_2~FF_brt_65 .SR_VALUE = 1'b0;
    defparam \RES[31]_2~FF_brt_65 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[31]_2~FF_brt_64  (.D(n5304), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[31]_2~FF_brt_64_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[31]_2~FF_brt_64 .CLK_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_64 .CE_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_64 .SR_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_64 .D_POLARITY = 1'b1;
    defparam \RES[31]_2~FF_brt_64 .SR_SYNC = 1'b1;
    defparam \RES[31]_2~FF_brt_64 .SR_VALUE = 1'b0;
    defparam \RES[31]_2~FF_brt_64 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[3]_2~FF_brt_121  (.D(n4949), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[3]_2~FF_brt_121_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[3]_2~FF_brt_121 .CLK_POLARITY = 1'b1;
    defparam \RES[3]_2~FF_brt_121 .CE_POLARITY = 1'b1;
    defparam \RES[3]_2~FF_brt_121 .SR_POLARITY = 1'b1;
    defparam \RES[3]_2~FF_brt_121 .D_POLARITY = 1'b1;
    defparam \RES[3]_2~FF_brt_121 .SR_SYNC = 1'b1;
    defparam \RES[3]_2~FF_brt_121 .SR_VALUE = 1'b0;
    defparam \RES[3]_2~FF_brt_121 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[29]_2~FF_brt_16_brt_62  (.D(n5283), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[29]_2~FF_brt_16_brt_62_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[29]_2~FF_brt_16_brt_62 .CLK_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_62 .CE_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_62 .SR_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_62 .D_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_62 .SR_SYNC = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_62 .SR_VALUE = 1'b0;
    defparam \RES[29]_2~FF_brt_16_brt_62 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[29]_2~FF_brt_16_brt_61  (.D(n5103), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[29]_2~FF_brt_16_brt_61_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[29]_2~FF_brt_16_brt_61 .CLK_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_61 .CE_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_61 .SR_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_61 .D_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_61 .SR_SYNC = 1'b1;
    defparam \RES[29]_2~FF_brt_16_brt_61 .SR_VALUE = 1'b0;
    defparam \RES[29]_2~FF_brt_16_brt_61 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_15_brt_59  (.D(n3445), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[28]_2~FF_brt_15_brt_59_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_15_brt_59 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_59 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_59 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_59 .D_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_59 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_59 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_15_brt_59 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_15_brt_58  (.D(n5275), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[28]_2~FF_brt_15_brt_58_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_15_brt_58 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_58 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_58 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_58 .D_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_58 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_58 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_15_brt_58 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_15_brt_57  (.D(n5276), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[28]_2~FF_brt_15_brt_57_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_15_brt_57 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_57 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_57 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_57 .D_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_57 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_15_brt_57 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_15_brt_57 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[27]_2~FF_brt_56  (.D(n5268), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[27]_2~FF_brt_56_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[27]_2~FF_brt_56 .CLK_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_56 .CE_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_56 .SR_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_56 .D_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_56 .SR_SYNC = 1'b1;
    defparam \RES[27]_2~FF_brt_56 .SR_VALUE = 1'b0;
    defparam \RES[27]_2~FF_brt_56 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[4]_2~FF_brt_123  (.D(n4964), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[4]_2~FF_brt_123_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[4]_2~FF_brt_123 .CLK_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_123 .CE_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_123 .SR_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_123 .D_POLARITY = 1'b0;
    defparam \RES[4]_2~FF_brt_123 .SR_SYNC = 1'b1;
    defparam \RES[4]_2~FF_brt_123 .SR_VALUE = 1'b0;
    defparam \RES[4]_2~FF_brt_123 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[27]_2~FF_brt_54  (.D(n5067), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[27]_2~FF_brt_54_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[27]_2~FF_brt_54 .CLK_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_54 .CE_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_54 .SR_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_54 .D_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_54 .SR_SYNC = 1'b1;
    defparam \RES[27]_2~FF_brt_54 .SR_VALUE = 1'b0;
    defparam \RES[27]_2~FF_brt_54 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[27]_2~FF_brt_53  (.D(n5075), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[27]_2~FF_brt_53_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[27]_2~FF_brt_53 .CLK_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_53 .CE_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_53 .SR_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_53 .D_POLARITY = 1'b1;
    defparam \RES[27]_2~FF_brt_53 .SR_SYNC = 1'b1;
    defparam \RES[27]_2~FF_brt_53 .SR_VALUE = 1'b0;
    defparam \RES[27]_2~FF_brt_53 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[4]_2~FF_brt_124  (.D(n4966), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[4]_2~FF_brt_124_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[4]_2~FF_brt_124 .CLK_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_124 .CE_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_124 .SR_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_124 .D_POLARITY = 1'b1;
    defparam \RES[4]_2~FF_brt_124 .SR_SYNC = 1'b1;
    defparam \RES[4]_2~FF_brt_124 .SR_VALUE = 1'b0;
    defparam \RES[4]_2~FF_brt_124 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[26]_2~FF_brt_10_brt_51  (.D(n5253), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[26]_2~FF_brt_10_brt_51_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[26]_2~FF_brt_10_brt_51 .CLK_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_51 .CE_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_51 .SR_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_51 .D_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_51 .SR_SYNC = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_51 .SR_VALUE = 1'b0;
    defparam \RES[26]_2~FF_brt_10_brt_51 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[26]_2~FF_brt_10_brt_50  (.D(n5249), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[26]_2~FF_brt_10_brt_50_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[26]_2~FF_brt_10_brt_50 .CLK_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_50 .CE_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_50 .SR_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_50 .D_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_50 .SR_SYNC = 1'b1;
    defparam \RES[26]_2~FF_brt_10_brt_50 .SR_VALUE = 1'b0;
    defparam \RES[26]_2~FF_brt_10_brt_50 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[5]_2~FF_brt_126  (.D(n4971), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[5]_2~FF_brt_126_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[5]_2~FF_brt_126 .CLK_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_126 .CE_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_126 .SR_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_126 .D_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_126 .SR_SYNC = 1'b1;
    defparam \RES[5]_2~FF_brt_126 .SR_VALUE = 1'b0;
    defparam \RES[5]_2~FF_brt_126 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_48  (.D(n3537), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[24]_2~FF_brt_48_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_48 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_48 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_48 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_48 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_48 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_48 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_48 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_47  (.D(n5225), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[24]_2~FF_brt_47_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_47 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_47 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_47 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_47 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_47 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_47 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_47 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[24]_2~FF_brt_46  (.D(n5224), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[24]_2~FF_brt_46_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[24]_2~FF_brt_46 .CLK_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_46 .CE_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_46 .SR_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_46 .D_POLARITY = 1'b1;
    defparam \RES[24]_2~FF_brt_46 .SR_SYNC = 1'b1;
    defparam \RES[24]_2~FF_brt_46 .SR_VALUE = 1'b0;
    defparam \RES[24]_2~FF_brt_46 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[5]_2~FF_brt_127  (.D(n4981), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[5]_2~FF_brt_127_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[5]_2~FF_brt_127 .CLK_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_127 .CE_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_127 .SR_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_127 .D_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_127 .SR_SYNC = 1'b1;
    defparam \RES[5]_2~FF_brt_127 .SR_VALUE = 1'b0;
    defparam \RES[5]_2~FF_brt_127 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[23]_2~FF_brt_44  (.D(n5213), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[23]_2~FF_brt_44_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[23]_2~FF_brt_44 .CLK_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_44 .CE_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_44 .SR_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_44 .D_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_44 .SR_SYNC = 1'b1;
    defparam \RES[23]_2~FF_brt_44 .SR_VALUE = 1'b0;
    defparam \RES[23]_2~FF_brt_44 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[23]_2~FF_brt_43  (.D(n5220), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[23]_2~FF_brt_43_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[23]_2~FF_brt_43 .CLK_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_43 .CE_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_43 .SR_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_43 .D_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_43 .SR_SYNC = 1'b1;
    defparam \RES[23]_2~FF_brt_43 .SR_VALUE = 1'b0;
    defparam \RES[23]_2~FF_brt_43 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[23]_2~FF_brt_42  (.D(n5218), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[23]_2~FF_brt_42_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[23]_2~FF_brt_42 .CLK_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_42 .CE_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_42 .SR_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_42 .D_POLARITY = 1'b1;
    defparam \RES[23]_2~FF_brt_42 .SR_SYNC = 1'b1;
    defparam \RES[23]_2~FF_brt_42 .SR_VALUE = 1'b0;
    defparam \RES[23]_2~FF_brt_42 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[5]_2~FF_brt_128  (.D(n4983), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[5]_2~FF_brt_128_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[5]_2~FF_brt_128 .CLK_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_128 .CE_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_128 .SR_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_128 .D_POLARITY = 1'b1;
    defparam \RES[5]_2~FF_brt_128 .SR_SYNC = 1'b1;
    defparam \RES[5]_2~FF_brt_128 .SR_VALUE = 1'b0;
    defparam \RES[5]_2~FF_brt_128 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[22]_2~FF_brt_39  (.D(n5212), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[22]_2~FF_brt_39_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[22]_2~FF_brt_39 .CLK_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_39 .CE_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_39 .SR_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_39 .D_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_39 .SR_SYNC = 1'b1;
    defparam \RES[22]_2~FF_brt_39 .SR_VALUE = 1'b0;
    defparam \RES[22]_2~FF_brt_39 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[22]_2~FF_brt_38  (.D(n5207), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[22]_2~FF_brt_38_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[22]_2~FF_brt_38 .CLK_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_38 .CE_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_38 .SR_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_38 .D_POLARITY = 1'b1;
    defparam \RES[22]_2~FF_brt_38 .SR_SYNC = 1'b1;
    defparam \RES[22]_2~FF_brt_38 .SR_VALUE = 1'b0;
    defparam \RES[22]_2~FF_brt_38 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[7]_2~FF_brt_20_brt_70_brt_132  (.D(n5017), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[7]_2~FF_brt_20_brt_70_brt_132_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_132 .CLK_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_132 .CE_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_132 .SR_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_132 .D_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_132 .SR_SYNC = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_132 .SR_VALUE = 1'b0;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_132 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_8_brt_36  (.D(\OPERATION[2] ), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[17]_2~FF_brt_8_brt_36_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_8_brt_36 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_36 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_36 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_36 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_36 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_36 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_8_brt_36 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_8_brt_35  (.D(n5145), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[17]_2~FF_brt_8_brt_35_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_8_brt_35 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_35 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_35 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_35 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_35 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_35 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_8_brt_35 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_8_brt_34  (.D(n4957), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[17]_2~FF_brt_8_brt_34_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_8_brt_34 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_34 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_34 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_34 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_34 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_8_brt_34 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_8_brt_34 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[7]_2~FF_brt_20_brt_70_brt_133  (.D(n5019), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[7]_2~FF_brt_20_brt_70_brt_133_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133 .CLK_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133 .CE_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133 .SR_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133 .D_POLARITY = 1'b0;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133 .SR_SYNC = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133 .SR_VALUE = 1'b0;
    defparam \RES[7]_2~FF_brt_20_brt_70_brt_133 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[16]_2~FF_brt_5_brt_32  (.D(n5135), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[16]_2~FF_brt_5_brt_32_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[16]_2~FF_brt_5_brt_32 .CLK_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_32 .CE_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_32 .SR_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_32 .D_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_32 .SR_SYNC = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_32 .SR_VALUE = 1'b0;
    defparam \RES[16]_2~FF_brt_5_brt_32 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[16]_2~FF_brt_5_brt_31  (.D(n5131), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[16]_2~FF_brt_5_brt_31_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[16]_2~FF_brt_5_brt_31 .CLK_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_31 .CE_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_31 .SR_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_31 .D_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_31 .SR_SYNC = 1'b1;
    defparam \RES[16]_2~FF_brt_5_brt_31 .SR_VALUE = 1'b0;
    defparam \RES[16]_2~FF_brt_5_brt_31 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[8]_2~FF_brt_21_brt_73_brt_134  (.D(n5033), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[8]_2~FF_brt_21_brt_73_brt_134_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[8]_2~FF_brt_21_brt_73_brt_134 .CLK_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_73_brt_134 .CE_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_73_brt_134 .SR_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_73_brt_134 .D_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_73_brt_134 .SR_SYNC = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_73_brt_134 .SR_VALUE = 1'b0;
    defparam \RES[8]_2~FF_brt_21_brt_73_brt_134 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[15]_2~FF_brt_29  (.D(n5123), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[15]_2~FF_brt_29_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[15]_2~FF_brt_29 .CLK_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_29 .CE_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_29 .SR_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_29 .D_POLARITY = 1'b0;
    defparam \RES[15]_2~FF_brt_29 .SR_SYNC = 1'b1;
    defparam \RES[15]_2~FF_brt_29 .SR_VALUE = 1'b0;
    defparam \RES[15]_2~FF_brt_29 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136  (.D(n1432), .CE(ceg_net408), 
           .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136 .D_POLARITY = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_136 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[10]_2~FF_brt_3_brt_27  (.D(n5053), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[10]_2~FF_brt_3_brt_27_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[10]_2~FF_brt_3_brt_27 .CLK_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_27 .CE_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_27 .SR_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_27 .D_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_27 .SR_SYNC = 1'b1;
    defparam \RES[10]_2~FF_brt_3_brt_27 .SR_VALUE = 1'b0;
    defparam \RES[10]_2~FF_brt_3_brt_27 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137  (.D(\OPERATION[1] ), 
           .CE(ceg_net408), .CLK(\CLK~O ), .SR(1'b0), .Q(\RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137 .D_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_26_brt_74_brt_137 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[9]_2~FF_brt_1_brt_25  (.D(n5046), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[9]_2~FF_brt_1_brt_25_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_1_brt_25 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_25 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_25 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_25 .D_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_25 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_1_brt_25 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_1_brt_25 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[29]_2~FF_brt_17  (.D(n5289), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[29]_2~FF_brt_17_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[29]_2~FF_brt_17 .CLK_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_17 .CE_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_17 .SR_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_17 .D_POLARITY = 1'b1;
    defparam \RES[29]_2~FF_brt_17 .SR_SYNC = 1'b1;
    defparam \RES[29]_2~FF_brt_17 .SR_VALUE = 1'b0;
    defparam \RES[29]_2~FF_brt_17 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[7]_2~FF_brt_20_brt_69  (.D(n5011), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[7]_2~FF_brt_20_brt_69_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[7]_2~FF_brt_20_brt_69 .CLK_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_69 .CE_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_69 .SR_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_69 .D_POLARITY = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_69 .SR_SYNC = 1'b1;
    defparam \RES[7]_2~FF_brt_20_brt_69 .SR_VALUE = 1'b0;
    defparam \RES[7]_2~FF_brt_20_brt_69 .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i30  (.I0(n2744), .I1(1'b1), .CI(1'b0), 
            .CO(n5924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i30 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i30 .I1_POLARITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_14  (.D(n3545), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[28]_2~FF_brt_14_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_14 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_14 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_14 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_14 .D_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_14 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_14 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_14 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[28]_2~FF_brt_13  (.D(n5271), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[28]_2~FF_brt_13_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[28]_2~FF_brt_13 .CLK_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_13 .CE_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_13 .SR_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_13 .D_POLARITY = 1'b1;
    defparam \RES[28]_2~FF_brt_13 .SR_SYNC = 1'b1;
    defparam \RES[28]_2~FF_brt_13 .SR_VALUE = 1'b0;
    defparam \RES[28]_2~FF_brt_13 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[26]_2~FF_brt_12  (.D(n5258), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[26]_2~FF_brt_12_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[26]_2~FF_brt_12 .CLK_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_12 .CE_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_12 .SR_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_12 .D_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_12 .SR_SYNC = 1'b1;
    defparam \RES[26]_2~FF_brt_12 .SR_VALUE = 1'b0;
    defparam \RES[26]_2~FF_brt_12 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[26]_2~FF_brt_11  (.D(n5248), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[26]_2~FF_brt_11_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[26]_2~FF_brt_11 .CLK_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_11 .CE_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_11 .SR_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_11 .D_POLARITY = 1'b1;
    defparam \RES[26]_2~FF_brt_11 .SR_SYNC = 1'b1;
    defparam \RES[26]_2~FF_brt_11 .SR_VALUE = 1'b0;
    defparam \RES[26]_2~FF_brt_11 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[8]_2~FF_brt_21_brt_72  (.D(n5032), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[8]_2~FF_brt_21_brt_72_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[8]_2~FF_brt_21_brt_72 .CLK_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_72 .CE_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_72 .SR_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_72 .D_POLARITY = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_72 .SR_SYNC = 1'b1;
    defparam \RES[8]_2~FF_brt_21_brt_72 .SR_VALUE = 1'b0;
    defparam \RES[8]_2~FF_brt_21_brt_72 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_9  (.D(n5155), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[17]_2~FF_brt_9_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_9 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_9 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_9 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_9 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_9 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_9 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_9 .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_184/add_2/i1  (.I0(1'b1), .I1(1'b1), .CI(1'b0), 
            .CO(n5921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(570)
    defparam \AUX_ADD_CI__sub_184/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_184/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_FF \RES[17]_2~FF_brt_7  (.D(n5152), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[17]_2~FF_brt_7_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[17]_2~FF_brt_7 .CLK_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_7 .CE_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_7 .SR_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_7 .D_POLARITY = 1'b1;
    defparam \RES[17]_2~FF_brt_7 .SR_SYNC = 1'b1;
    defparam \RES[17]_2~FF_brt_7 .SR_VALUE = 1'b0;
    defparam \RES[17]_2~FF_brt_7 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[16]_2~FF_brt_6  (.D(n5141), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[16]_2~FF_brt_6_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[16]_2~FF_brt_6 .CLK_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_6 .CE_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_6 .SR_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_6 .D_POLARITY = 1'b1;
    defparam \RES[16]_2~FF_brt_6 .SR_SYNC = 1'b1;
    defparam \RES[16]_2~FF_brt_6 .SR_VALUE = 1'b0;
    defparam \RES[16]_2~FF_brt_6 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[12]_2~FF_brt_77  (.D(n5083), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[12]_2~FF_brt_77_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[12]_2~FF_brt_77 .CLK_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_77 .CE_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_77 .SR_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_77 .D_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_77 .SR_SYNC = 1'b1;
    defparam \RES[12]_2~FF_brt_77 .SR_VALUE = 1'b0;
    defparam \RES[12]_2~FF_brt_77 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[10]_2~FF_brt_4  (.D(n5063), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[10]_2~FF_brt_4_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[10]_2~FF_brt_4 .CLK_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_4 .CE_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_4 .SR_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_4 .D_POLARITY = 1'b1;
    defparam \RES[10]_2~FF_brt_4 .SR_SYNC = 1'b1;
    defparam \RES[10]_2~FF_brt_4 .SR_VALUE = 1'b0;
    defparam \RES[10]_2~FF_brt_4 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[12]_2~FF_brt_79  (.D(n5093), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[12]_2~FF_brt_79_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[12]_2~FF_brt_79 .CLK_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_79 .CE_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_79 .SR_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_79 .D_POLARITY = 1'b1;
    defparam \RES[12]_2~FF_brt_79 .SR_SYNC = 1'b1;
    defparam \RES[12]_2~FF_brt_79 .SR_VALUE = 1'b0;
    defparam \RES[12]_2~FF_brt_79 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[15]_2~FF_brt_30_brt_80  (.D(n5121), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[15]_2~FF_brt_30_brt_80_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[15]_2~FF_brt_30_brt_80 .CLK_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_80 .CE_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_80 .SR_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_80 .D_POLARITY = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_80 .SR_SYNC = 1'b1;
    defparam \RES[15]_2~FF_brt_30_brt_80 .SR_VALUE = 1'b0;
    defparam \RES[15]_2~FF_brt_30_brt_80 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RES[9]_2~FF_brt_0  (.D(n5041), .CE(ceg_net408), .CLK(\CLK~O ), 
           .SR(1'b0), .Q(\RES[9]_2~FF_brt_0_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Efinity\2022.1\project\New_RiscV\RISC_V_core.vhd(593)
    defparam \RES[9]_2~FF_brt_0 .CLK_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_0 .CE_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_0 .SR_POLARITY = 1'b1;
    defparam \RES[9]_2~FF_brt_0 .D_POLARITY = 1'b0;
    defparam \RES[9]_2~FF_brt_0 .SR_SYNC = 1'b1;
    defparam \RES[9]_2~FF_brt_0 .SR_VALUE = 1'b0;
    defparam \RES[9]_2~FF_brt_0 .SR_SYNC_PRIORITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bb0b1060_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bb0b1060_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bb0b1060_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bb0b1060_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_bb0b1060_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_bb0b1060_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__4_4_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__4_4_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__5_5_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__5_5_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__5_5_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__5_5_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__4_4_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bb0b1060__2_2_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bb0b1060_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_bb0b1060_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bb0b1060_4
// module not written out since it is a black box. 
//

